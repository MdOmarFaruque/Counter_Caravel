magic
tech sky130A
magscale 1 2
timestamp 1707334428
<< nwell >>
rect 1066 47045 18898 47366
rect 1066 45957 18898 46523
rect 1066 44869 18898 45435
rect 1066 43781 18898 44347
rect 1066 42693 18898 43259
rect 1066 41605 18898 42171
rect 1066 40517 18898 41083
rect 1066 39429 18898 39995
rect 1066 38341 18898 38907
rect 1066 37253 18898 37819
rect 1066 36165 18898 36731
rect 1066 35077 18898 35643
rect 1066 33989 18898 34555
rect 1066 32901 18898 33467
rect 1066 31813 18898 32379
rect 1066 30725 18898 31291
rect 1066 29637 18898 30203
rect 1066 28549 18898 29115
rect 1066 27461 18898 28027
rect 1066 26373 18898 26939
rect 1066 25285 18898 25851
rect 1066 24197 18898 24763
rect 1066 23109 18898 23675
rect 1066 22021 18898 22587
rect 1066 20933 18898 21499
rect 1066 19845 18898 20411
rect 1066 18757 18898 19323
rect 1066 17669 18898 18235
rect 1066 16581 18898 17147
rect 1066 15493 18898 16059
rect 1066 14405 18898 14971
rect 1066 13317 18898 13883
rect 1066 12229 18898 12795
rect 1066 11141 18898 11707
rect 1066 10053 18898 10619
rect 1066 8965 18898 9531
rect 1066 7877 18898 8443
rect 1066 6789 18898 7355
rect 1066 5701 18898 6267
rect 1066 4613 18898 5179
rect 1066 3525 18898 4091
rect 1066 2437 18898 3003
<< obsli1 >>
rect 1104 2159 18860 47345
<< obsm1 >>
rect 1104 2128 19019 47376
<< metal2 >>
rect 4986 0 5042 800
rect 14922 0 14978 800
<< obsm2 >>
rect 3169 856 19013 47365
rect 3169 800 4930 856
rect 5098 800 14866 856
rect 15034 800 19013 856
<< metal3 >>
rect 19200 46792 20000 46912
rect 19200 40536 20000 40656
rect 19200 34280 20000 34400
rect 19200 28024 20000 28144
rect 19200 21768 20000 21888
rect 19200 15512 20000 15632
rect 19200 9256 20000 9376
rect 19200 3000 20000 3120
<< obsm3 >>
rect 3165 46992 19626 47361
rect 3165 46712 19120 46992
rect 3165 40736 19626 46712
rect 3165 40456 19120 40736
rect 3165 34480 19626 40456
rect 3165 34200 19120 34480
rect 3165 28224 19626 34200
rect 3165 27944 19120 28224
rect 3165 21968 19626 27944
rect 3165 21688 19120 21968
rect 3165 15712 19626 21688
rect 3165 15432 19120 15712
rect 3165 9456 19626 15432
rect 3165 9176 19120 9456
rect 3165 3200 19626 9176
rect 3165 2920 19120 3200
rect 3165 2143 19626 2920
<< metal4 >>
rect 3163 2128 3483 47376
rect 5382 2128 5702 47376
rect 7602 2128 7922 47376
rect 9821 2128 10141 47376
rect 12041 2128 12361 47376
rect 14260 2128 14580 47376
rect 16480 2128 16800 47376
rect 18699 2128 19019 47376
<< labels >>
rlabel metal3 s 19200 9256 20000 9376 6 io_oeb[0]
port 1 nsew signal output
rlabel metal3 s 19200 21768 20000 21888 6 io_oeb[1]
port 2 nsew signal output
rlabel metal3 s 19200 34280 20000 34400 6 io_oeb[2]
port 3 nsew signal output
rlabel metal3 s 19200 46792 20000 46912 6 io_oeb[3]
port 4 nsew signal output
rlabel metal3 s 19200 3000 20000 3120 6 io_out[0]
port 5 nsew signal output
rlabel metal3 s 19200 15512 20000 15632 6 io_out[1]
port 6 nsew signal output
rlabel metal3 s 19200 28024 20000 28144 6 io_out[2]
port 7 nsew signal output
rlabel metal3 s 19200 40536 20000 40656 6 io_out[3]
port 8 nsew signal output
rlabel metal4 s 3163 2128 3483 47376 6 vccd1
port 9 nsew power bidirectional
rlabel metal4 s 7602 2128 7922 47376 6 vccd1
port 9 nsew power bidirectional
rlabel metal4 s 12041 2128 12361 47376 6 vccd1
port 9 nsew power bidirectional
rlabel metal4 s 16480 2128 16800 47376 6 vccd1
port 9 nsew power bidirectional
rlabel metal4 s 5382 2128 5702 47376 6 vssd1
port 10 nsew ground bidirectional
rlabel metal4 s 9821 2128 10141 47376 6 vssd1
port 10 nsew ground bidirectional
rlabel metal4 s 14260 2128 14580 47376 6 vssd1
port 10 nsew ground bidirectional
rlabel metal4 s 18699 2128 19019 47376 6 vssd1
port 10 nsew ground bidirectional
rlabel metal2 s 4986 0 5042 800 6 wb_clk_i
port 11 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wb_rst_i
port 12 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 682744
string GDS_FILE /home/engtech/Desktop/Openlane_v2/counter_v2/openlane/user_proj_example/runs/24_02_07_13_32/results/signoff/user_proj_example.magic.gds
string GDS_START 130470
<< end >>

