VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 46.280 100.000 46.880 ;
    END
  END io_oeb[0]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 108.840 100.000 109.440 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 171.400 100.000 172.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 233.960 100.000 234.560 ;
    END
  END io_oeb[3]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 15.000 100.000 15.600 ;
    END
  END io_out[0]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.560 100.000 78.160 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 140.120 100.000 140.720 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 96.000 202.680 100.000 203.280 ;
    END
  END io_out[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.815 10.640 17.415 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.010 10.640 39.610 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.205 10.640 61.805 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.400 10.640 84.000 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 26.910 10.640 28.510 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.105 10.640 50.705 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.300 10.640 72.900 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.495 10.640 95.095 236.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wb_rst_i
  OBS
      LAYER nwell ;
        RECT 5.330 235.225 94.490 236.830 ;
        RECT 5.330 229.785 94.490 232.615 ;
        RECT 5.330 224.345 94.490 227.175 ;
        RECT 5.330 218.905 94.490 221.735 ;
        RECT 5.330 213.465 94.490 216.295 ;
        RECT 5.330 208.025 94.490 210.855 ;
        RECT 5.330 202.585 94.490 205.415 ;
        RECT 5.330 197.145 94.490 199.975 ;
        RECT 5.330 191.705 94.490 194.535 ;
        RECT 5.330 186.265 94.490 189.095 ;
        RECT 5.330 180.825 94.490 183.655 ;
        RECT 5.330 175.385 94.490 178.215 ;
        RECT 5.330 169.945 94.490 172.775 ;
        RECT 5.330 164.505 94.490 167.335 ;
        RECT 5.330 159.065 94.490 161.895 ;
        RECT 5.330 153.625 94.490 156.455 ;
        RECT 5.330 148.185 94.490 151.015 ;
        RECT 5.330 142.745 94.490 145.575 ;
        RECT 5.330 137.305 94.490 140.135 ;
        RECT 5.330 131.865 94.490 134.695 ;
        RECT 5.330 126.425 94.490 129.255 ;
        RECT 5.330 120.985 94.490 123.815 ;
        RECT 5.330 115.545 94.490 118.375 ;
        RECT 5.330 110.105 94.490 112.935 ;
        RECT 5.330 104.665 94.490 107.495 ;
        RECT 5.330 99.225 94.490 102.055 ;
        RECT 5.330 93.785 94.490 96.615 ;
        RECT 5.330 88.345 94.490 91.175 ;
        RECT 5.330 82.905 94.490 85.735 ;
        RECT 5.330 77.465 94.490 80.295 ;
        RECT 5.330 72.025 94.490 74.855 ;
        RECT 5.330 66.585 94.490 69.415 ;
        RECT 5.330 61.145 94.490 63.975 ;
        RECT 5.330 55.705 94.490 58.535 ;
        RECT 5.330 50.265 94.490 53.095 ;
        RECT 5.330 44.825 94.490 47.655 ;
        RECT 5.330 39.385 94.490 42.215 ;
        RECT 5.330 33.945 94.490 36.775 ;
        RECT 5.330 28.505 94.490 31.335 ;
        RECT 5.330 23.065 94.490 25.895 ;
        RECT 5.330 17.625 94.490 20.455 ;
        RECT 5.330 12.185 94.490 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 94.300 236.725 ;
      LAYER met1 ;
        RECT 5.520 10.640 95.095 236.880 ;
      LAYER met2 ;
        RECT 15.845 4.280 95.065 236.825 ;
        RECT 15.845 4.000 24.650 4.280 ;
        RECT 25.490 4.000 74.330 4.280 ;
        RECT 75.170 4.000 95.065 4.280 ;
      LAYER met3 ;
        RECT 15.825 234.960 98.130 236.805 ;
        RECT 15.825 233.560 95.600 234.960 ;
        RECT 15.825 203.680 98.130 233.560 ;
        RECT 15.825 202.280 95.600 203.680 ;
        RECT 15.825 172.400 98.130 202.280 ;
        RECT 15.825 171.000 95.600 172.400 ;
        RECT 15.825 141.120 98.130 171.000 ;
        RECT 15.825 139.720 95.600 141.120 ;
        RECT 15.825 109.840 98.130 139.720 ;
        RECT 15.825 108.440 95.600 109.840 ;
        RECT 15.825 78.560 98.130 108.440 ;
        RECT 15.825 77.160 95.600 78.560 ;
        RECT 15.825 47.280 98.130 77.160 ;
        RECT 15.825 45.880 95.600 47.280 ;
        RECT 15.825 16.000 98.130 45.880 ;
        RECT 15.825 14.600 95.600 16.000 ;
        RECT 15.825 10.715 98.130 14.600 ;
  END
END user_proj_example
END LIBRARY

