magic
tech sky130A
magscale 1 2
timestamp 1707334427
<< viali >>
rect 18521 47209 18555 47243
rect 18337 41089 18371 41123
rect 17877 41021 17911 41055
rect 18429 40341 18463 40375
rect 18521 34357 18555 34391
rect 17141 28509 17175 28543
rect 18337 28441 18371 28475
rect 17049 28373 17083 28407
rect 18521 22185 18555 22219
rect 17141 16065 17175 16099
rect 18337 15997 18371 16031
rect 18521 9333 18555 9367
rect 18429 8585 18463 8619
rect 15945 8517 15979 8551
rect 15761 8449 15795 8483
rect 16037 8449 16071 8483
rect 15761 8313 15795 8347
rect 16037 7973 16071 8007
rect 17417 7905 17451 7939
rect 18429 7905 18463 7939
rect 15853 7837 15887 7871
rect 16773 7837 16807 7871
rect 17693 7837 17727 7871
rect 17785 7837 17819 7871
rect 15669 7701 15703 7735
rect 16129 7701 16163 7735
rect 17417 7701 17451 7735
rect 17601 7701 17635 7735
rect 17877 7701 17911 7735
rect 14933 7497 14967 7531
rect 18337 7497 18371 7531
rect 16057 7361 16091 7395
rect 16957 7361 16991 7395
rect 17224 7361 17258 7395
rect 16313 7293 16347 7327
rect 17417 6953 17451 6987
rect 17601 6953 17635 6987
rect 15669 6817 15703 6851
rect 16221 6817 16255 6851
rect 16405 6817 16439 6851
rect 16589 6817 16623 6851
rect 16773 6817 16807 6851
rect 17877 6817 17911 6851
rect 17969 6817 18003 6851
rect 18153 6817 18187 6851
rect 15393 6749 15427 6783
rect 15577 6749 15611 6783
rect 16681 6749 16715 6783
rect 16865 6749 16899 6783
rect 17049 6749 17083 6783
rect 18061 6749 18095 6783
rect 15485 6613 15519 6647
rect 17417 6613 17451 6647
rect 17693 6613 17727 6647
rect 16129 5865 16163 5899
rect 17417 5593 17451 5627
rect 16129 5321 16163 5355
rect 15945 5253 15979 5287
rect 16221 5185 16255 5219
rect 16681 5185 16715 5219
rect 15945 4981 15979 5015
rect 17969 4981 18003 5015
rect 15761 4573 15795 4607
rect 17325 4573 17359 4607
rect 17601 4573 17635 4607
rect 16028 4505 16062 4539
rect 17141 4437 17175 4471
rect 15945 4233 15979 4267
rect 16129 4097 16163 4131
rect 16313 4097 16347 4131
rect 16405 4097 16439 4131
rect 17325 4097 17359 4131
rect 18337 4029 18371 4063
rect 17509 3689 17543 3723
rect 18245 3621 18279 3655
rect 18061 3553 18095 3587
rect 17417 3485 17451 3519
rect 18429 3417 18463 3451
rect 16129 3349 16163 3383
rect 18061 3145 18095 3179
rect 16405 3077 16439 3111
rect 16926 3077 16960 3111
rect 16313 3009 16347 3043
rect 16497 3009 16531 3043
rect 16681 2941 16715 2975
rect 15209 2601 15243 2635
rect 18521 2601 18555 2635
rect 17877 2465 17911 2499
rect 15025 2397 15059 2431
<< metal1 >>
rect 1104 47354 18860 47376
rect 1104 47302 3169 47354
rect 3221 47302 3233 47354
rect 3285 47302 3297 47354
rect 3349 47302 3361 47354
rect 3413 47302 3425 47354
rect 3477 47302 7608 47354
rect 7660 47302 7672 47354
rect 7724 47302 7736 47354
rect 7788 47302 7800 47354
rect 7852 47302 7864 47354
rect 7916 47302 12047 47354
rect 12099 47302 12111 47354
rect 12163 47302 12175 47354
rect 12227 47302 12239 47354
rect 12291 47302 12303 47354
rect 12355 47302 16486 47354
rect 16538 47302 16550 47354
rect 16602 47302 16614 47354
rect 16666 47302 16678 47354
rect 16730 47302 16742 47354
rect 16794 47302 18860 47354
rect 1104 47280 18860 47302
rect 18506 47200 18512 47252
rect 18564 47200 18570 47252
rect 1104 46810 19019 46832
rect 1104 46758 5388 46810
rect 5440 46758 5452 46810
rect 5504 46758 5516 46810
rect 5568 46758 5580 46810
rect 5632 46758 5644 46810
rect 5696 46758 9827 46810
rect 9879 46758 9891 46810
rect 9943 46758 9955 46810
rect 10007 46758 10019 46810
rect 10071 46758 10083 46810
rect 10135 46758 14266 46810
rect 14318 46758 14330 46810
rect 14382 46758 14394 46810
rect 14446 46758 14458 46810
rect 14510 46758 14522 46810
rect 14574 46758 18705 46810
rect 18757 46758 18769 46810
rect 18821 46758 18833 46810
rect 18885 46758 18897 46810
rect 18949 46758 18961 46810
rect 19013 46758 19019 46810
rect 1104 46736 19019 46758
rect 1104 46266 18860 46288
rect 1104 46214 3169 46266
rect 3221 46214 3233 46266
rect 3285 46214 3297 46266
rect 3349 46214 3361 46266
rect 3413 46214 3425 46266
rect 3477 46214 7608 46266
rect 7660 46214 7672 46266
rect 7724 46214 7736 46266
rect 7788 46214 7800 46266
rect 7852 46214 7864 46266
rect 7916 46214 12047 46266
rect 12099 46214 12111 46266
rect 12163 46214 12175 46266
rect 12227 46214 12239 46266
rect 12291 46214 12303 46266
rect 12355 46214 16486 46266
rect 16538 46214 16550 46266
rect 16602 46214 16614 46266
rect 16666 46214 16678 46266
rect 16730 46214 16742 46266
rect 16794 46214 18860 46266
rect 1104 46192 18860 46214
rect 1104 45722 19019 45744
rect 1104 45670 5388 45722
rect 5440 45670 5452 45722
rect 5504 45670 5516 45722
rect 5568 45670 5580 45722
rect 5632 45670 5644 45722
rect 5696 45670 9827 45722
rect 9879 45670 9891 45722
rect 9943 45670 9955 45722
rect 10007 45670 10019 45722
rect 10071 45670 10083 45722
rect 10135 45670 14266 45722
rect 14318 45670 14330 45722
rect 14382 45670 14394 45722
rect 14446 45670 14458 45722
rect 14510 45670 14522 45722
rect 14574 45670 18705 45722
rect 18757 45670 18769 45722
rect 18821 45670 18833 45722
rect 18885 45670 18897 45722
rect 18949 45670 18961 45722
rect 19013 45670 19019 45722
rect 1104 45648 19019 45670
rect 1104 45178 18860 45200
rect 1104 45126 3169 45178
rect 3221 45126 3233 45178
rect 3285 45126 3297 45178
rect 3349 45126 3361 45178
rect 3413 45126 3425 45178
rect 3477 45126 7608 45178
rect 7660 45126 7672 45178
rect 7724 45126 7736 45178
rect 7788 45126 7800 45178
rect 7852 45126 7864 45178
rect 7916 45126 12047 45178
rect 12099 45126 12111 45178
rect 12163 45126 12175 45178
rect 12227 45126 12239 45178
rect 12291 45126 12303 45178
rect 12355 45126 16486 45178
rect 16538 45126 16550 45178
rect 16602 45126 16614 45178
rect 16666 45126 16678 45178
rect 16730 45126 16742 45178
rect 16794 45126 18860 45178
rect 1104 45104 18860 45126
rect 1104 44634 19019 44656
rect 1104 44582 5388 44634
rect 5440 44582 5452 44634
rect 5504 44582 5516 44634
rect 5568 44582 5580 44634
rect 5632 44582 5644 44634
rect 5696 44582 9827 44634
rect 9879 44582 9891 44634
rect 9943 44582 9955 44634
rect 10007 44582 10019 44634
rect 10071 44582 10083 44634
rect 10135 44582 14266 44634
rect 14318 44582 14330 44634
rect 14382 44582 14394 44634
rect 14446 44582 14458 44634
rect 14510 44582 14522 44634
rect 14574 44582 18705 44634
rect 18757 44582 18769 44634
rect 18821 44582 18833 44634
rect 18885 44582 18897 44634
rect 18949 44582 18961 44634
rect 19013 44582 19019 44634
rect 1104 44560 19019 44582
rect 1104 44090 18860 44112
rect 1104 44038 3169 44090
rect 3221 44038 3233 44090
rect 3285 44038 3297 44090
rect 3349 44038 3361 44090
rect 3413 44038 3425 44090
rect 3477 44038 7608 44090
rect 7660 44038 7672 44090
rect 7724 44038 7736 44090
rect 7788 44038 7800 44090
rect 7852 44038 7864 44090
rect 7916 44038 12047 44090
rect 12099 44038 12111 44090
rect 12163 44038 12175 44090
rect 12227 44038 12239 44090
rect 12291 44038 12303 44090
rect 12355 44038 16486 44090
rect 16538 44038 16550 44090
rect 16602 44038 16614 44090
rect 16666 44038 16678 44090
rect 16730 44038 16742 44090
rect 16794 44038 18860 44090
rect 1104 44016 18860 44038
rect 1104 43546 19019 43568
rect 1104 43494 5388 43546
rect 5440 43494 5452 43546
rect 5504 43494 5516 43546
rect 5568 43494 5580 43546
rect 5632 43494 5644 43546
rect 5696 43494 9827 43546
rect 9879 43494 9891 43546
rect 9943 43494 9955 43546
rect 10007 43494 10019 43546
rect 10071 43494 10083 43546
rect 10135 43494 14266 43546
rect 14318 43494 14330 43546
rect 14382 43494 14394 43546
rect 14446 43494 14458 43546
rect 14510 43494 14522 43546
rect 14574 43494 18705 43546
rect 18757 43494 18769 43546
rect 18821 43494 18833 43546
rect 18885 43494 18897 43546
rect 18949 43494 18961 43546
rect 19013 43494 19019 43546
rect 1104 43472 19019 43494
rect 1104 43002 18860 43024
rect 1104 42950 3169 43002
rect 3221 42950 3233 43002
rect 3285 42950 3297 43002
rect 3349 42950 3361 43002
rect 3413 42950 3425 43002
rect 3477 42950 7608 43002
rect 7660 42950 7672 43002
rect 7724 42950 7736 43002
rect 7788 42950 7800 43002
rect 7852 42950 7864 43002
rect 7916 42950 12047 43002
rect 12099 42950 12111 43002
rect 12163 42950 12175 43002
rect 12227 42950 12239 43002
rect 12291 42950 12303 43002
rect 12355 42950 16486 43002
rect 16538 42950 16550 43002
rect 16602 42950 16614 43002
rect 16666 42950 16678 43002
rect 16730 42950 16742 43002
rect 16794 42950 18860 43002
rect 1104 42928 18860 42950
rect 1104 42458 19019 42480
rect 1104 42406 5388 42458
rect 5440 42406 5452 42458
rect 5504 42406 5516 42458
rect 5568 42406 5580 42458
rect 5632 42406 5644 42458
rect 5696 42406 9827 42458
rect 9879 42406 9891 42458
rect 9943 42406 9955 42458
rect 10007 42406 10019 42458
rect 10071 42406 10083 42458
rect 10135 42406 14266 42458
rect 14318 42406 14330 42458
rect 14382 42406 14394 42458
rect 14446 42406 14458 42458
rect 14510 42406 14522 42458
rect 14574 42406 18705 42458
rect 18757 42406 18769 42458
rect 18821 42406 18833 42458
rect 18885 42406 18897 42458
rect 18949 42406 18961 42458
rect 19013 42406 19019 42458
rect 1104 42384 19019 42406
rect 1104 41914 18860 41936
rect 1104 41862 3169 41914
rect 3221 41862 3233 41914
rect 3285 41862 3297 41914
rect 3349 41862 3361 41914
rect 3413 41862 3425 41914
rect 3477 41862 7608 41914
rect 7660 41862 7672 41914
rect 7724 41862 7736 41914
rect 7788 41862 7800 41914
rect 7852 41862 7864 41914
rect 7916 41862 12047 41914
rect 12099 41862 12111 41914
rect 12163 41862 12175 41914
rect 12227 41862 12239 41914
rect 12291 41862 12303 41914
rect 12355 41862 16486 41914
rect 16538 41862 16550 41914
rect 16602 41862 16614 41914
rect 16666 41862 16678 41914
rect 16730 41862 16742 41914
rect 16794 41862 18860 41914
rect 1104 41840 18860 41862
rect 1104 41370 19019 41392
rect 1104 41318 5388 41370
rect 5440 41318 5452 41370
rect 5504 41318 5516 41370
rect 5568 41318 5580 41370
rect 5632 41318 5644 41370
rect 5696 41318 9827 41370
rect 9879 41318 9891 41370
rect 9943 41318 9955 41370
rect 10007 41318 10019 41370
rect 10071 41318 10083 41370
rect 10135 41318 14266 41370
rect 14318 41318 14330 41370
rect 14382 41318 14394 41370
rect 14446 41318 14458 41370
rect 14510 41318 14522 41370
rect 14574 41318 18705 41370
rect 18757 41318 18769 41370
rect 18821 41318 18833 41370
rect 18885 41318 18897 41370
rect 18949 41318 18961 41370
rect 19013 41318 19019 41370
rect 1104 41296 19019 41318
rect 18322 41080 18328 41132
rect 18380 41080 18386 41132
rect 17865 41055 17923 41061
rect 17865 41021 17877 41055
rect 17911 41052 17923 41055
rect 18046 41052 18052 41064
rect 17911 41024 18052 41052
rect 17911 41021 17923 41024
rect 17865 41015 17923 41021
rect 18046 41012 18052 41024
rect 18104 41012 18110 41064
rect 1104 40826 18860 40848
rect 1104 40774 3169 40826
rect 3221 40774 3233 40826
rect 3285 40774 3297 40826
rect 3349 40774 3361 40826
rect 3413 40774 3425 40826
rect 3477 40774 7608 40826
rect 7660 40774 7672 40826
rect 7724 40774 7736 40826
rect 7788 40774 7800 40826
rect 7852 40774 7864 40826
rect 7916 40774 12047 40826
rect 12099 40774 12111 40826
rect 12163 40774 12175 40826
rect 12227 40774 12239 40826
rect 12291 40774 12303 40826
rect 12355 40774 16486 40826
rect 16538 40774 16550 40826
rect 16602 40774 16614 40826
rect 16666 40774 16678 40826
rect 16730 40774 16742 40826
rect 16794 40774 18860 40826
rect 1104 40752 18860 40774
rect 18322 40332 18328 40384
rect 18380 40372 18386 40384
rect 18417 40375 18475 40381
rect 18417 40372 18429 40375
rect 18380 40344 18429 40372
rect 18380 40332 18386 40344
rect 18417 40341 18429 40344
rect 18463 40341 18475 40375
rect 18417 40335 18475 40341
rect 1104 40282 19019 40304
rect 1104 40230 5388 40282
rect 5440 40230 5452 40282
rect 5504 40230 5516 40282
rect 5568 40230 5580 40282
rect 5632 40230 5644 40282
rect 5696 40230 9827 40282
rect 9879 40230 9891 40282
rect 9943 40230 9955 40282
rect 10007 40230 10019 40282
rect 10071 40230 10083 40282
rect 10135 40230 14266 40282
rect 14318 40230 14330 40282
rect 14382 40230 14394 40282
rect 14446 40230 14458 40282
rect 14510 40230 14522 40282
rect 14574 40230 18705 40282
rect 18757 40230 18769 40282
rect 18821 40230 18833 40282
rect 18885 40230 18897 40282
rect 18949 40230 18961 40282
rect 19013 40230 19019 40282
rect 1104 40208 19019 40230
rect 1104 39738 18860 39760
rect 1104 39686 3169 39738
rect 3221 39686 3233 39738
rect 3285 39686 3297 39738
rect 3349 39686 3361 39738
rect 3413 39686 3425 39738
rect 3477 39686 7608 39738
rect 7660 39686 7672 39738
rect 7724 39686 7736 39738
rect 7788 39686 7800 39738
rect 7852 39686 7864 39738
rect 7916 39686 12047 39738
rect 12099 39686 12111 39738
rect 12163 39686 12175 39738
rect 12227 39686 12239 39738
rect 12291 39686 12303 39738
rect 12355 39686 16486 39738
rect 16538 39686 16550 39738
rect 16602 39686 16614 39738
rect 16666 39686 16678 39738
rect 16730 39686 16742 39738
rect 16794 39686 18860 39738
rect 1104 39664 18860 39686
rect 1104 39194 19019 39216
rect 1104 39142 5388 39194
rect 5440 39142 5452 39194
rect 5504 39142 5516 39194
rect 5568 39142 5580 39194
rect 5632 39142 5644 39194
rect 5696 39142 9827 39194
rect 9879 39142 9891 39194
rect 9943 39142 9955 39194
rect 10007 39142 10019 39194
rect 10071 39142 10083 39194
rect 10135 39142 14266 39194
rect 14318 39142 14330 39194
rect 14382 39142 14394 39194
rect 14446 39142 14458 39194
rect 14510 39142 14522 39194
rect 14574 39142 18705 39194
rect 18757 39142 18769 39194
rect 18821 39142 18833 39194
rect 18885 39142 18897 39194
rect 18949 39142 18961 39194
rect 19013 39142 19019 39194
rect 1104 39120 19019 39142
rect 1104 38650 18860 38672
rect 1104 38598 3169 38650
rect 3221 38598 3233 38650
rect 3285 38598 3297 38650
rect 3349 38598 3361 38650
rect 3413 38598 3425 38650
rect 3477 38598 7608 38650
rect 7660 38598 7672 38650
rect 7724 38598 7736 38650
rect 7788 38598 7800 38650
rect 7852 38598 7864 38650
rect 7916 38598 12047 38650
rect 12099 38598 12111 38650
rect 12163 38598 12175 38650
rect 12227 38598 12239 38650
rect 12291 38598 12303 38650
rect 12355 38598 16486 38650
rect 16538 38598 16550 38650
rect 16602 38598 16614 38650
rect 16666 38598 16678 38650
rect 16730 38598 16742 38650
rect 16794 38598 18860 38650
rect 1104 38576 18860 38598
rect 1104 38106 19019 38128
rect 1104 38054 5388 38106
rect 5440 38054 5452 38106
rect 5504 38054 5516 38106
rect 5568 38054 5580 38106
rect 5632 38054 5644 38106
rect 5696 38054 9827 38106
rect 9879 38054 9891 38106
rect 9943 38054 9955 38106
rect 10007 38054 10019 38106
rect 10071 38054 10083 38106
rect 10135 38054 14266 38106
rect 14318 38054 14330 38106
rect 14382 38054 14394 38106
rect 14446 38054 14458 38106
rect 14510 38054 14522 38106
rect 14574 38054 18705 38106
rect 18757 38054 18769 38106
rect 18821 38054 18833 38106
rect 18885 38054 18897 38106
rect 18949 38054 18961 38106
rect 19013 38054 19019 38106
rect 1104 38032 19019 38054
rect 1104 37562 18860 37584
rect 1104 37510 3169 37562
rect 3221 37510 3233 37562
rect 3285 37510 3297 37562
rect 3349 37510 3361 37562
rect 3413 37510 3425 37562
rect 3477 37510 7608 37562
rect 7660 37510 7672 37562
rect 7724 37510 7736 37562
rect 7788 37510 7800 37562
rect 7852 37510 7864 37562
rect 7916 37510 12047 37562
rect 12099 37510 12111 37562
rect 12163 37510 12175 37562
rect 12227 37510 12239 37562
rect 12291 37510 12303 37562
rect 12355 37510 16486 37562
rect 16538 37510 16550 37562
rect 16602 37510 16614 37562
rect 16666 37510 16678 37562
rect 16730 37510 16742 37562
rect 16794 37510 18860 37562
rect 1104 37488 18860 37510
rect 1104 37018 19019 37040
rect 1104 36966 5388 37018
rect 5440 36966 5452 37018
rect 5504 36966 5516 37018
rect 5568 36966 5580 37018
rect 5632 36966 5644 37018
rect 5696 36966 9827 37018
rect 9879 36966 9891 37018
rect 9943 36966 9955 37018
rect 10007 36966 10019 37018
rect 10071 36966 10083 37018
rect 10135 36966 14266 37018
rect 14318 36966 14330 37018
rect 14382 36966 14394 37018
rect 14446 36966 14458 37018
rect 14510 36966 14522 37018
rect 14574 36966 18705 37018
rect 18757 36966 18769 37018
rect 18821 36966 18833 37018
rect 18885 36966 18897 37018
rect 18949 36966 18961 37018
rect 19013 36966 19019 37018
rect 1104 36944 19019 36966
rect 1104 36474 18860 36496
rect 1104 36422 3169 36474
rect 3221 36422 3233 36474
rect 3285 36422 3297 36474
rect 3349 36422 3361 36474
rect 3413 36422 3425 36474
rect 3477 36422 7608 36474
rect 7660 36422 7672 36474
rect 7724 36422 7736 36474
rect 7788 36422 7800 36474
rect 7852 36422 7864 36474
rect 7916 36422 12047 36474
rect 12099 36422 12111 36474
rect 12163 36422 12175 36474
rect 12227 36422 12239 36474
rect 12291 36422 12303 36474
rect 12355 36422 16486 36474
rect 16538 36422 16550 36474
rect 16602 36422 16614 36474
rect 16666 36422 16678 36474
rect 16730 36422 16742 36474
rect 16794 36422 18860 36474
rect 1104 36400 18860 36422
rect 1104 35930 19019 35952
rect 1104 35878 5388 35930
rect 5440 35878 5452 35930
rect 5504 35878 5516 35930
rect 5568 35878 5580 35930
rect 5632 35878 5644 35930
rect 5696 35878 9827 35930
rect 9879 35878 9891 35930
rect 9943 35878 9955 35930
rect 10007 35878 10019 35930
rect 10071 35878 10083 35930
rect 10135 35878 14266 35930
rect 14318 35878 14330 35930
rect 14382 35878 14394 35930
rect 14446 35878 14458 35930
rect 14510 35878 14522 35930
rect 14574 35878 18705 35930
rect 18757 35878 18769 35930
rect 18821 35878 18833 35930
rect 18885 35878 18897 35930
rect 18949 35878 18961 35930
rect 19013 35878 19019 35930
rect 1104 35856 19019 35878
rect 1104 35386 18860 35408
rect 1104 35334 3169 35386
rect 3221 35334 3233 35386
rect 3285 35334 3297 35386
rect 3349 35334 3361 35386
rect 3413 35334 3425 35386
rect 3477 35334 7608 35386
rect 7660 35334 7672 35386
rect 7724 35334 7736 35386
rect 7788 35334 7800 35386
rect 7852 35334 7864 35386
rect 7916 35334 12047 35386
rect 12099 35334 12111 35386
rect 12163 35334 12175 35386
rect 12227 35334 12239 35386
rect 12291 35334 12303 35386
rect 12355 35334 16486 35386
rect 16538 35334 16550 35386
rect 16602 35334 16614 35386
rect 16666 35334 16678 35386
rect 16730 35334 16742 35386
rect 16794 35334 18860 35386
rect 1104 35312 18860 35334
rect 1104 34842 19019 34864
rect 1104 34790 5388 34842
rect 5440 34790 5452 34842
rect 5504 34790 5516 34842
rect 5568 34790 5580 34842
rect 5632 34790 5644 34842
rect 5696 34790 9827 34842
rect 9879 34790 9891 34842
rect 9943 34790 9955 34842
rect 10007 34790 10019 34842
rect 10071 34790 10083 34842
rect 10135 34790 14266 34842
rect 14318 34790 14330 34842
rect 14382 34790 14394 34842
rect 14446 34790 14458 34842
rect 14510 34790 14522 34842
rect 14574 34790 18705 34842
rect 18757 34790 18769 34842
rect 18821 34790 18833 34842
rect 18885 34790 18897 34842
rect 18949 34790 18961 34842
rect 19013 34790 19019 34842
rect 1104 34768 19019 34790
rect 18506 34348 18512 34400
rect 18564 34348 18570 34400
rect 1104 34298 18860 34320
rect 1104 34246 3169 34298
rect 3221 34246 3233 34298
rect 3285 34246 3297 34298
rect 3349 34246 3361 34298
rect 3413 34246 3425 34298
rect 3477 34246 7608 34298
rect 7660 34246 7672 34298
rect 7724 34246 7736 34298
rect 7788 34246 7800 34298
rect 7852 34246 7864 34298
rect 7916 34246 12047 34298
rect 12099 34246 12111 34298
rect 12163 34246 12175 34298
rect 12227 34246 12239 34298
rect 12291 34246 12303 34298
rect 12355 34246 16486 34298
rect 16538 34246 16550 34298
rect 16602 34246 16614 34298
rect 16666 34246 16678 34298
rect 16730 34246 16742 34298
rect 16794 34246 18860 34298
rect 1104 34224 18860 34246
rect 1104 33754 19019 33776
rect 1104 33702 5388 33754
rect 5440 33702 5452 33754
rect 5504 33702 5516 33754
rect 5568 33702 5580 33754
rect 5632 33702 5644 33754
rect 5696 33702 9827 33754
rect 9879 33702 9891 33754
rect 9943 33702 9955 33754
rect 10007 33702 10019 33754
rect 10071 33702 10083 33754
rect 10135 33702 14266 33754
rect 14318 33702 14330 33754
rect 14382 33702 14394 33754
rect 14446 33702 14458 33754
rect 14510 33702 14522 33754
rect 14574 33702 18705 33754
rect 18757 33702 18769 33754
rect 18821 33702 18833 33754
rect 18885 33702 18897 33754
rect 18949 33702 18961 33754
rect 19013 33702 19019 33754
rect 1104 33680 19019 33702
rect 1104 33210 18860 33232
rect 1104 33158 3169 33210
rect 3221 33158 3233 33210
rect 3285 33158 3297 33210
rect 3349 33158 3361 33210
rect 3413 33158 3425 33210
rect 3477 33158 7608 33210
rect 7660 33158 7672 33210
rect 7724 33158 7736 33210
rect 7788 33158 7800 33210
rect 7852 33158 7864 33210
rect 7916 33158 12047 33210
rect 12099 33158 12111 33210
rect 12163 33158 12175 33210
rect 12227 33158 12239 33210
rect 12291 33158 12303 33210
rect 12355 33158 16486 33210
rect 16538 33158 16550 33210
rect 16602 33158 16614 33210
rect 16666 33158 16678 33210
rect 16730 33158 16742 33210
rect 16794 33158 18860 33210
rect 1104 33136 18860 33158
rect 1104 32666 19019 32688
rect 1104 32614 5388 32666
rect 5440 32614 5452 32666
rect 5504 32614 5516 32666
rect 5568 32614 5580 32666
rect 5632 32614 5644 32666
rect 5696 32614 9827 32666
rect 9879 32614 9891 32666
rect 9943 32614 9955 32666
rect 10007 32614 10019 32666
rect 10071 32614 10083 32666
rect 10135 32614 14266 32666
rect 14318 32614 14330 32666
rect 14382 32614 14394 32666
rect 14446 32614 14458 32666
rect 14510 32614 14522 32666
rect 14574 32614 18705 32666
rect 18757 32614 18769 32666
rect 18821 32614 18833 32666
rect 18885 32614 18897 32666
rect 18949 32614 18961 32666
rect 19013 32614 19019 32666
rect 1104 32592 19019 32614
rect 1104 32122 18860 32144
rect 1104 32070 3169 32122
rect 3221 32070 3233 32122
rect 3285 32070 3297 32122
rect 3349 32070 3361 32122
rect 3413 32070 3425 32122
rect 3477 32070 7608 32122
rect 7660 32070 7672 32122
rect 7724 32070 7736 32122
rect 7788 32070 7800 32122
rect 7852 32070 7864 32122
rect 7916 32070 12047 32122
rect 12099 32070 12111 32122
rect 12163 32070 12175 32122
rect 12227 32070 12239 32122
rect 12291 32070 12303 32122
rect 12355 32070 16486 32122
rect 16538 32070 16550 32122
rect 16602 32070 16614 32122
rect 16666 32070 16678 32122
rect 16730 32070 16742 32122
rect 16794 32070 18860 32122
rect 1104 32048 18860 32070
rect 1104 31578 19019 31600
rect 1104 31526 5388 31578
rect 5440 31526 5452 31578
rect 5504 31526 5516 31578
rect 5568 31526 5580 31578
rect 5632 31526 5644 31578
rect 5696 31526 9827 31578
rect 9879 31526 9891 31578
rect 9943 31526 9955 31578
rect 10007 31526 10019 31578
rect 10071 31526 10083 31578
rect 10135 31526 14266 31578
rect 14318 31526 14330 31578
rect 14382 31526 14394 31578
rect 14446 31526 14458 31578
rect 14510 31526 14522 31578
rect 14574 31526 18705 31578
rect 18757 31526 18769 31578
rect 18821 31526 18833 31578
rect 18885 31526 18897 31578
rect 18949 31526 18961 31578
rect 19013 31526 19019 31578
rect 1104 31504 19019 31526
rect 1104 31034 18860 31056
rect 1104 30982 3169 31034
rect 3221 30982 3233 31034
rect 3285 30982 3297 31034
rect 3349 30982 3361 31034
rect 3413 30982 3425 31034
rect 3477 30982 7608 31034
rect 7660 30982 7672 31034
rect 7724 30982 7736 31034
rect 7788 30982 7800 31034
rect 7852 30982 7864 31034
rect 7916 30982 12047 31034
rect 12099 30982 12111 31034
rect 12163 30982 12175 31034
rect 12227 30982 12239 31034
rect 12291 30982 12303 31034
rect 12355 30982 16486 31034
rect 16538 30982 16550 31034
rect 16602 30982 16614 31034
rect 16666 30982 16678 31034
rect 16730 30982 16742 31034
rect 16794 30982 18860 31034
rect 1104 30960 18860 30982
rect 1104 30490 19019 30512
rect 1104 30438 5388 30490
rect 5440 30438 5452 30490
rect 5504 30438 5516 30490
rect 5568 30438 5580 30490
rect 5632 30438 5644 30490
rect 5696 30438 9827 30490
rect 9879 30438 9891 30490
rect 9943 30438 9955 30490
rect 10007 30438 10019 30490
rect 10071 30438 10083 30490
rect 10135 30438 14266 30490
rect 14318 30438 14330 30490
rect 14382 30438 14394 30490
rect 14446 30438 14458 30490
rect 14510 30438 14522 30490
rect 14574 30438 18705 30490
rect 18757 30438 18769 30490
rect 18821 30438 18833 30490
rect 18885 30438 18897 30490
rect 18949 30438 18961 30490
rect 19013 30438 19019 30490
rect 1104 30416 19019 30438
rect 1104 29946 18860 29968
rect 1104 29894 3169 29946
rect 3221 29894 3233 29946
rect 3285 29894 3297 29946
rect 3349 29894 3361 29946
rect 3413 29894 3425 29946
rect 3477 29894 7608 29946
rect 7660 29894 7672 29946
rect 7724 29894 7736 29946
rect 7788 29894 7800 29946
rect 7852 29894 7864 29946
rect 7916 29894 12047 29946
rect 12099 29894 12111 29946
rect 12163 29894 12175 29946
rect 12227 29894 12239 29946
rect 12291 29894 12303 29946
rect 12355 29894 16486 29946
rect 16538 29894 16550 29946
rect 16602 29894 16614 29946
rect 16666 29894 16678 29946
rect 16730 29894 16742 29946
rect 16794 29894 18860 29946
rect 1104 29872 18860 29894
rect 1104 29402 19019 29424
rect 1104 29350 5388 29402
rect 5440 29350 5452 29402
rect 5504 29350 5516 29402
rect 5568 29350 5580 29402
rect 5632 29350 5644 29402
rect 5696 29350 9827 29402
rect 9879 29350 9891 29402
rect 9943 29350 9955 29402
rect 10007 29350 10019 29402
rect 10071 29350 10083 29402
rect 10135 29350 14266 29402
rect 14318 29350 14330 29402
rect 14382 29350 14394 29402
rect 14446 29350 14458 29402
rect 14510 29350 14522 29402
rect 14574 29350 18705 29402
rect 18757 29350 18769 29402
rect 18821 29350 18833 29402
rect 18885 29350 18897 29402
rect 18949 29350 18961 29402
rect 19013 29350 19019 29402
rect 1104 29328 19019 29350
rect 1104 28858 18860 28880
rect 1104 28806 3169 28858
rect 3221 28806 3233 28858
rect 3285 28806 3297 28858
rect 3349 28806 3361 28858
rect 3413 28806 3425 28858
rect 3477 28806 7608 28858
rect 7660 28806 7672 28858
rect 7724 28806 7736 28858
rect 7788 28806 7800 28858
rect 7852 28806 7864 28858
rect 7916 28806 12047 28858
rect 12099 28806 12111 28858
rect 12163 28806 12175 28858
rect 12227 28806 12239 28858
rect 12291 28806 12303 28858
rect 12355 28806 16486 28858
rect 16538 28806 16550 28858
rect 16602 28806 16614 28858
rect 16666 28806 16678 28858
rect 16730 28806 16742 28858
rect 16794 28806 18860 28858
rect 1104 28784 18860 28806
rect 17129 28543 17187 28549
rect 17129 28540 17141 28543
rect 17052 28512 17141 28540
rect 17052 28416 17080 28512
rect 17129 28509 17141 28512
rect 17175 28509 17187 28543
rect 17129 28503 17187 28509
rect 18325 28475 18383 28481
rect 18325 28441 18337 28475
rect 18371 28472 18383 28475
rect 18598 28472 18604 28484
rect 18371 28444 18604 28472
rect 18371 28441 18383 28444
rect 18325 28435 18383 28441
rect 18598 28432 18604 28444
rect 18656 28432 18662 28484
rect 17034 28364 17040 28416
rect 17092 28364 17098 28416
rect 1104 28314 19019 28336
rect 1104 28262 5388 28314
rect 5440 28262 5452 28314
rect 5504 28262 5516 28314
rect 5568 28262 5580 28314
rect 5632 28262 5644 28314
rect 5696 28262 9827 28314
rect 9879 28262 9891 28314
rect 9943 28262 9955 28314
rect 10007 28262 10019 28314
rect 10071 28262 10083 28314
rect 10135 28262 14266 28314
rect 14318 28262 14330 28314
rect 14382 28262 14394 28314
rect 14446 28262 14458 28314
rect 14510 28262 14522 28314
rect 14574 28262 18705 28314
rect 18757 28262 18769 28314
rect 18821 28262 18833 28314
rect 18885 28262 18897 28314
rect 18949 28262 18961 28314
rect 19013 28262 19019 28314
rect 1104 28240 19019 28262
rect 1104 27770 18860 27792
rect 1104 27718 3169 27770
rect 3221 27718 3233 27770
rect 3285 27718 3297 27770
rect 3349 27718 3361 27770
rect 3413 27718 3425 27770
rect 3477 27718 7608 27770
rect 7660 27718 7672 27770
rect 7724 27718 7736 27770
rect 7788 27718 7800 27770
rect 7852 27718 7864 27770
rect 7916 27718 12047 27770
rect 12099 27718 12111 27770
rect 12163 27718 12175 27770
rect 12227 27718 12239 27770
rect 12291 27718 12303 27770
rect 12355 27718 16486 27770
rect 16538 27718 16550 27770
rect 16602 27718 16614 27770
rect 16666 27718 16678 27770
rect 16730 27718 16742 27770
rect 16794 27718 18860 27770
rect 1104 27696 18860 27718
rect 1104 27226 19019 27248
rect 1104 27174 5388 27226
rect 5440 27174 5452 27226
rect 5504 27174 5516 27226
rect 5568 27174 5580 27226
rect 5632 27174 5644 27226
rect 5696 27174 9827 27226
rect 9879 27174 9891 27226
rect 9943 27174 9955 27226
rect 10007 27174 10019 27226
rect 10071 27174 10083 27226
rect 10135 27174 14266 27226
rect 14318 27174 14330 27226
rect 14382 27174 14394 27226
rect 14446 27174 14458 27226
rect 14510 27174 14522 27226
rect 14574 27174 18705 27226
rect 18757 27174 18769 27226
rect 18821 27174 18833 27226
rect 18885 27174 18897 27226
rect 18949 27174 18961 27226
rect 19013 27174 19019 27226
rect 1104 27152 19019 27174
rect 1104 26682 18860 26704
rect 1104 26630 3169 26682
rect 3221 26630 3233 26682
rect 3285 26630 3297 26682
rect 3349 26630 3361 26682
rect 3413 26630 3425 26682
rect 3477 26630 7608 26682
rect 7660 26630 7672 26682
rect 7724 26630 7736 26682
rect 7788 26630 7800 26682
rect 7852 26630 7864 26682
rect 7916 26630 12047 26682
rect 12099 26630 12111 26682
rect 12163 26630 12175 26682
rect 12227 26630 12239 26682
rect 12291 26630 12303 26682
rect 12355 26630 16486 26682
rect 16538 26630 16550 26682
rect 16602 26630 16614 26682
rect 16666 26630 16678 26682
rect 16730 26630 16742 26682
rect 16794 26630 18860 26682
rect 1104 26608 18860 26630
rect 1104 26138 19019 26160
rect 1104 26086 5388 26138
rect 5440 26086 5452 26138
rect 5504 26086 5516 26138
rect 5568 26086 5580 26138
rect 5632 26086 5644 26138
rect 5696 26086 9827 26138
rect 9879 26086 9891 26138
rect 9943 26086 9955 26138
rect 10007 26086 10019 26138
rect 10071 26086 10083 26138
rect 10135 26086 14266 26138
rect 14318 26086 14330 26138
rect 14382 26086 14394 26138
rect 14446 26086 14458 26138
rect 14510 26086 14522 26138
rect 14574 26086 18705 26138
rect 18757 26086 18769 26138
rect 18821 26086 18833 26138
rect 18885 26086 18897 26138
rect 18949 26086 18961 26138
rect 19013 26086 19019 26138
rect 1104 26064 19019 26086
rect 1104 25594 18860 25616
rect 1104 25542 3169 25594
rect 3221 25542 3233 25594
rect 3285 25542 3297 25594
rect 3349 25542 3361 25594
rect 3413 25542 3425 25594
rect 3477 25542 7608 25594
rect 7660 25542 7672 25594
rect 7724 25542 7736 25594
rect 7788 25542 7800 25594
rect 7852 25542 7864 25594
rect 7916 25542 12047 25594
rect 12099 25542 12111 25594
rect 12163 25542 12175 25594
rect 12227 25542 12239 25594
rect 12291 25542 12303 25594
rect 12355 25542 16486 25594
rect 16538 25542 16550 25594
rect 16602 25542 16614 25594
rect 16666 25542 16678 25594
rect 16730 25542 16742 25594
rect 16794 25542 18860 25594
rect 1104 25520 18860 25542
rect 1104 25050 19019 25072
rect 1104 24998 5388 25050
rect 5440 24998 5452 25050
rect 5504 24998 5516 25050
rect 5568 24998 5580 25050
rect 5632 24998 5644 25050
rect 5696 24998 9827 25050
rect 9879 24998 9891 25050
rect 9943 24998 9955 25050
rect 10007 24998 10019 25050
rect 10071 24998 10083 25050
rect 10135 24998 14266 25050
rect 14318 24998 14330 25050
rect 14382 24998 14394 25050
rect 14446 24998 14458 25050
rect 14510 24998 14522 25050
rect 14574 24998 18705 25050
rect 18757 24998 18769 25050
rect 18821 24998 18833 25050
rect 18885 24998 18897 25050
rect 18949 24998 18961 25050
rect 19013 24998 19019 25050
rect 1104 24976 19019 24998
rect 1104 24506 18860 24528
rect 1104 24454 3169 24506
rect 3221 24454 3233 24506
rect 3285 24454 3297 24506
rect 3349 24454 3361 24506
rect 3413 24454 3425 24506
rect 3477 24454 7608 24506
rect 7660 24454 7672 24506
rect 7724 24454 7736 24506
rect 7788 24454 7800 24506
rect 7852 24454 7864 24506
rect 7916 24454 12047 24506
rect 12099 24454 12111 24506
rect 12163 24454 12175 24506
rect 12227 24454 12239 24506
rect 12291 24454 12303 24506
rect 12355 24454 16486 24506
rect 16538 24454 16550 24506
rect 16602 24454 16614 24506
rect 16666 24454 16678 24506
rect 16730 24454 16742 24506
rect 16794 24454 18860 24506
rect 1104 24432 18860 24454
rect 1104 23962 19019 23984
rect 1104 23910 5388 23962
rect 5440 23910 5452 23962
rect 5504 23910 5516 23962
rect 5568 23910 5580 23962
rect 5632 23910 5644 23962
rect 5696 23910 9827 23962
rect 9879 23910 9891 23962
rect 9943 23910 9955 23962
rect 10007 23910 10019 23962
rect 10071 23910 10083 23962
rect 10135 23910 14266 23962
rect 14318 23910 14330 23962
rect 14382 23910 14394 23962
rect 14446 23910 14458 23962
rect 14510 23910 14522 23962
rect 14574 23910 18705 23962
rect 18757 23910 18769 23962
rect 18821 23910 18833 23962
rect 18885 23910 18897 23962
rect 18949 23910 18961 23962
rect 19013 23910 19019 23962
rect 1104 23888 19019 23910
rect 1104 23418 18860 23440
rect 1104 23366 3169 23418
rect 3221 23366 3233 23418
rect 3285 23366 3297 23418
rect 3349 23366 3361 23418
rect 3413 23366 3425 23418
rect 3477 23366 7608 23418
rect 7660 23366 7672 23418
rect 7724 23366 7736 23418
rect 7788 23366 7800 23418
rect 7852 23366 7864 23418
rect 7916 23366 12047 23418
rect 12099 23366 12111 23418
rect 12163 23366 12175 23418
rect 12227 23366 12239 23418
rect 12291 23366 12303 23418
rect 12355 23366 16486 23418
rect 16538 23366 16550 23418
rect 16602 23366 16614 23418
rect 16666 23366 16678 23418
rect 16730 23366 16742 23418
rect 16794 23366 18860 23418
rect 1104 23344 18860 23366
rect 1104 22874 19019 22896
rect 1104 22822 5388 22874
rect 5440 22822 5452 22874
rect 5504 22822 5516 22874
rect 5568 22822 5580 22874
rect 5632 22822 5644 22874
rect 5696 22822 9827 22874
rect 9879 22822 9891 22874
rect 9943 22822 9955 22874
rect 10007 22822 10019 22874
rect 10071 22822 10083 22874
rect 10135 22822 14266 22874
rect 14318 22822 14330 22874
rect 14382 22822 14394 22874
rect 14446 22822 14458 22874
rect 14510 22822 14522 22874
rect 14574 22822 18705 22874
rect 18757 22822 18769 22874
rect 18821 22822 18833 22874
rect 18885 22822 18897 22874
rect 18949 22822 18961 22874
rect 19013 22822 19019 22874
rect 1104 22800 19019 22822
rect 1104 22330 18860 22352
rect 1104 22278 3169 22330
rect 3221 22278 3233 22330
rect 3285 22278 3297 22330
rect 3349 22278 3361 22330
rect 3413 22278 3425 22330
rect 3477 22278 7608 22330
rect 7660 22278 7672 22330
rect 7724 22278 7736 22330
rect 7788 22278 7800 22330
rect 7852 22278 7864 22330
rect 7916 22278 12047 22330
rect 12099 22278 12111 22330
rect 12163 22278 12175 22330
rect 12227 22278 12239 22330
rect 12291 22278 12303 22330
rect 12355 22278 16486 22330
rect 16538 22278 16550 22330
rect 16602 22278 16614 22330
rect 16666 22278 16678 22330
rect 16730 22278 16742 22330
rect 16794 22278 18860 22330
rect 1104 22256 18860 22278
rect 18506 22176 18512 22228
rect 18564 22176 18570 22228
rect 1104 21786 19019 21808
rect 1104 21734 5388 21786
rect 5440 21734 5452 21786
rect 5504 21734 5516 21786
rect 5568 21734 5580 21786
rect 5632 21734 5644 21786
rect 5696 21734 9827 21786
rect 9879 21734 9891 21786
rect 9943 21734 9955 21786
rect 10007 21734 10019 21786
rect 10071 21734 10083 21786
rect 10135 21734 14266 21786
rect 14318 21734 14330 21786
rect 14382 21734 14394 21786
rect 14446 21734 14458 21786
rect 14510 21734 14522 21786
rect 14574 21734 18705 21786
rect 18757 21734 18769 21786
rect 18821 21734 18833 21786
rect 18885 21734 18897 21786
rect 18949 21734 18961 21786
rect 19013 21734 19019 21786
rect 1104 21712 19019 21734
rect 1104 21242 18860 21264
rect 1104 21190 3169 21242
rect 3221 21190 3233 21242
rect 3285 21190 3297 21242
rect 3349 21190 3361 21242
rect 3413 21190 3425 21242
rect 3477 21190 7608 21242
rect 7660 21190 7672 21242
rect 7724 21190 7736 21242
rect 7788 21190 7800 21242
rect 7852 21190 7864 21242
rect 7916 21190 12047 21242
rect 12099 21190 12111 21242
rect 12163 21190 12175 21242
rect 12227 21190 12239 21242
rect 12291 21190 12303 21242
rect 12355 21190 16486 21242
rect 16538 21190 16550 21242
rect 16602 21190 16614 21242
rect 16666 21190 16678 21242
rect 16730 21190 16742 21242
rect 16794 21190 18860 21242
rect 1104 21168 18860 21190
rect 1104 20698 19019 20720
rect 1104 20646 5388 20698
rect 5440 20646 5452 20698
rect 5504 20646 5516 20698
rect 5568 20646 5580 20698
rect 5632 20646 5644 20698
rect 5696 20646 9827 20698
rect 9879 20646 9891 20698
rect 9943 20646 9955 20698
rect 10007 20646 10019 20698
rect 10071 20646 10083 20698
rect 10135 20646 14266 20698
rect 14318 20646 14330 20698
rect 14382 20646 14394 20698
rect 14446 20646 14458 20698
rect 14510 20646 14522 20698
rect 14574 20646 18705 20698
rect 18757 20646 18769 20698
rect 18821 20646 18833 20698
rect 18885 20646 18897 20698
rect 18949 20646 18961 20698
rect 19013 20646 19019 20698
rect 1104 20624 19019 20646
rect 1104 20154 18860 20176
rect 1104 20102 3169 20154
rect 3221 20102 3233 20154
rect 3285 20102 3297 20154
rect 3349 20102 3361 20154
rect 3413 20102 3425 20154
rect 3477 20102 7608 20154
rect 7660 20102 7672 20154
rect 7724 20102 7736 20154
rect 7788 20102 7800 20154
rect 7852 20102 7864 20154
rect 7916 20102 12047 20154
rect 12099 20102 12111 20154
rect 12163 20102 12175 20154
rect 12227 20102 12239 20154
rect 12291 20102 12303 20154
rect 12355 20102 16486 20154
rect 16538 20102 16550 20154
rect 16602 20102 16614 20154
rect 16666 20102 16678 20154
rect 16730 20102 16742 20154
rect 16794 20102 18860 20154
rect 1104 20080 18860 20102
rect 1104 19610 19019 19632
rect 1104 19558 5388 19610
rect 5440 19558 5452 19610
rect 5504 19558 5516 19610
rect 5568 19558 5580 19610
rect 5632 19558 5644 19610
rect 5696 19558 9827 19610
rect 9879 19558 9891 19610
rect 9943 19558 9955 19610
rect 10007 19558 10019 19610
rect 10071 19558 10083 19610
rect 10135 19558 14266 19610
rect 14318 19558 14330 19610
rect 14382 19558 14394 19610
rect 14446 19558 14458 19610
rect 14510 19558 14522 19610
rect 14574 19558 18705 19610
rect 18757 19558 18769 19610
rect 18821 19558 18833 19610
rect 18885 19558 18897 19610
rect 18949 19558 18961 19610
rect 19013 19558 19019 19610
rect 1104 19536 19019 19558
rect 1104 19066 18860 19088
rect 1104 19014 3169 19066
rect 3221 19014 3233 19066
rect 3285 19014 3297 19066
rect 3349 19014 3361 19066
rect 3413 19014 3425 19066
rect 3477 19014 7608 19066
rect 7660 19014 7672 19066
rect 7724 19014 7736 19066
rect 7788 19014 7800 19066
rect 7852 19014 7864 19066
rect 7916 19014 12047 19066
rect 12099 19014 12111 19066
rect 12163 19014 12175 19066
rect 12227 19014 12239 19066
rect 12291 19014 12303 19066
rect 12355 19014 16486 19066
rect 16538 19014 16550 19066
rect 16602 19014 16614 19066
rect 16666 19014 16678 19066
rect 16730 19014 16742 19066
rect 16794 19014 18860 19066
rect 1104 18992 18860 19014
rect 1104 18522 19019 18544
rect 1104 18470 5388 18522
rect 5440 18470 5452 18522
rect 5504 18470 5516 18522
rect 5568 18470 5580 18522
rect 5632 18470 5644 18522
rect 5696 18470 9827 18522
rect 9879 18470 9891 18522
rect 9943 18470 9955 18522
rect 10007 18470 10019 18522
rect 10071 18470 10083 18522
rect 10135 18470 14266 18522
rect 14318 18470 14330 18522
rect 14382 18470 14394 18522
rect 14446 18470 14458 18522
rect 14510 18470 14522 18522
rect 14574 18470 18705 18522
rect 18757 18470 18769 18522
rect 18821 18470 18833 18522
rect 18885 18470 18897 18522
rect 18949 18470 18961 18522
rect 19013 18470 19019 18522
rect 1104 18448 19019 18470
rect 1104 17978 18860 18000
rect 1104 17926 3169 17978
rect 3221 17926 3233 17978
rect 3285 17926 3297 17978
rect 3349 17926 3361 17978
rect 3413 17926 3425 17978
rect 3477 17926 7608 17978
rect 7660 17926 7672 17978
rect 7724 17926 7736 17978
rect 7788 17926 7800 17978
rect 7852 17926 7864 17978
rect 7916 17926 12047 17978
rect 12099 17926 12111 17978
rect 12163 17926 12175 17978
rect 12227 17926 12239 17978
rect 12291 17926 12303 17978
rect 12355 17926 16486 17978
rect 16538 17926 16550 17978
rect 16602 17926 16614 17978
rect 16666 17926 16678 17978
rect 16730 17926 16742 17978
rect 16794 17926 18860 17978
rect 1104 17904 18860 17926
rect 1104 17434 19019 17456
rect 1104 17382 5388 17434
rect 5440 17382 5452 17434
rect 5504 17382 5516 17434
rect 5568 17382 5580 17434
rect 5632 17382 5644 17434
rect 5696 17382 9827 17434
rect 9879 17382 9891 17434
rect 9943 17382 9955 17434
rect 10007 17382 10019 17434
rect 10071 17382 10083 17434
rect 10135 17382 14266 17434
rect 14318 17382 14330 17434
rect 14382 17382 14394 17434
rect 14446 17382 14458 17434
rect 14510 17382 14522 17434
rect 14574 17382 18705 17434
rect 18757 17382 18769 17434
rect 18821 17382 18833 17434
rect 18885 17382 18897 17434
rect 18949 17382 18961 17434
rect 19013 17382 19019 17434
rect 1104 17360 19019 17382
rect 1104 16890 18860 16912
rect 1104 16838 3169 16890
rect 3221 16838 3233 16890
rect 3285 16838 3297 16890
rect 3349 16838 3361 16890
rect 3413 16838 3425 16890
rect 3477 16838 7608 16890
rect 7660 16838 7672 16890
rect 7724 16838 7736 16890
rect 7788 16838 7800 16890
rect 7852 16838 7864 16890
rect 7916 16838 12047 16890
rect 12099 16838 12111 16890
rect 12163 16838 12175 16890
rect 12227 16838 12239 16890
rect 12291 16838 12303 16890
rect 12355 16838 16486 16890
rect 16538 16838 16550 16890
rect 16602 16838 16614 16890
rect 16666 16838 16678 16890
rect 16730 16838 16742 16890
rect 16794 16838 18860 16890
rect 1104 16816 18860 16838
rect 1104 16346 19019 16368
rect 1104 16294 5388 16346
rect 5440 16294 5452 16346
rect 5504 16294 5516 16346
rect 5568 16294 5580 16346
rect 5632 16294 5644 16346
rect 5696 16294 9827 16346
rect 9879 16294 9891 16346
rect 9943 16294 9955 16346
rect 10007 16294 10019 16346
rect 10071 16294 10083 16346
rect 10135 16294 14266 16346
rect 14318 16294 14330 16346
rect 14382 16294 14394 16346
rect 14446 16294 14458 16346
rect 14510 16294 14522 16346
rect 14574 16294 18705 16346
rect 18757 16294 18769 16346
rect 18821 16294 18833 16346
rect 18885 16294 18897 16346
rect 18949 16294 18961 16346
rect 19013 16294 19019 16346
rect 1104 16272 19019 16294
rect 17126 16056 17132 16108
rect 17184 16056 17190 16108
rect 18322 15988 18328 16040
rect 18380 15988 18386 16040
rect 1104 15802 18860 15824
rect 1104 15750 3169 15802
rect 3221 15750 3233 15802
rect 3285 15750 3297 15802
rect 3349 15750 3361 15802
rect 3413 15750 3425 15802
rect 3477 15750 7608 15802
rect 7660 15750 7672 15802
rect 7724 15750 7736 15802
rect 7788 15750 7800 15802
rect 7852 15750 7864 15802
rect 7916 15750 12047 15802
rect 12099 15750 12111 15802
rect 12163 15750 12175 15802
rect 12227 15750 12239 15802
rect 12291 15750 12303 15802
rect 12355 15750 16486 15802
rect 16538 15750 16550 15802
rect 16602 15750 16614 15802
rect 16666 15750 16678 15802
rect 16730 15750 16742 15802
rect 16794 15750 18860 15802
rect 1104 15728 18860 15750
rect 1104 15258 19019 15280
rect 1104 15206 5388 15258
rect 5440 15206 5452 15258
rect 5504 15206 5516 15258
rect 5568 15206 5580 15258
rect 5632 15206 5644 15258
rect 5696 15206 9827 15258
rect 9879 15206 9891 15258
rect 9943 15206 9955 15258
rect 10007 15206 10019 15258
rect 10071 15206 10083 15258
rect 10135 15206 14266 15258
rect 14318 15206 14330 15258
rect 14382 15206 14394 15258
rect 14446 15206 14458 15258
rect 14510 15206 14522 15258
rect 14574 15206 18705 15258
rect 18757 15206 18769 15258
rect 18821 15206 18833 15258
rect 18885 15206 18897 15258
rect 18949 15206 18961 15258
rect 19013 15206 19019 15258
rect 1104 15184 19019 15206
rect 1104 14714 18860 14736
rect 1104 14662 3169 14714
rect 3221 14662 3233 14714
rect 3285 14662 3297 14714
rect 3349 14662 3361 14714
rect 3413 14662 3425 14714
rect 3477 14662 7608 14714
rect 7660 14662 7672 14714
rect 7724 14662 7736 14714
rect 7788 14662 7800 14714
rect 7852 14662 7864 14714
rect 7916 14662 12047 14714
rect 12099 14662 12111 14714
rect 12163 14662 12175 14714
rect 12227 14662 12239 14714
rect 12291 14662 12303 14714
rect 12355 14662 16486 14714
rect 16538 14662 16550 14714
rect 16602 14662 16614 14714
rect 16666 14662 16678 14714
rect 16730 14662 16742 14714
rect 16794 14662 18860 14714
rect 1104 14640 18860 14662
rect 1104 14170 19019 14192
rect 1104 14118 5388 14170
rect 5440 14118 5452 14170
rect 5504 14118 5516 14170
rect 5568 14118 5580 14170
rect 5632 14118 5644 14170
rect 5696 14118 9827 14170
rect 9879 14118 9891 14170
rect 9943 14118 9955 14170
rect 10007 14118 10019 14170
rect 10071 14118 10083 14170
rect 10135 14118 14266 14170
rect 14318 14118 14330 14170
rect 14382 14118 14394 14170
rect 14446 14118 14458 14170
rect 14510 14118 14522 14170
rect 14574 14118 18705 14170
rect 18757 14118 18769 14170
rect 18821 14118 18833 14170
rect 18885 14118 18897 14170
rect 18949 14118 18961 14170
rect 19013 14118 19019 14170
rect 1104 14096 19019 14118
rect 1104 13626 18860 13648
rect 1104 13574 3169 13626
rect 3221 13574 3233 13626
rect 3285 13574 3297 13626
rect 3349 13574 3361 13626
rect 3413 13574 3425 13626
rect 3477 13574 7608 13626
rect 7660 13574 7672 13626
rect 7724 13574 7736 13626
rect 7788 13574 7800 13626
rect 7852 13574 7864 13626
rect 7916 13574 12047 13626
rect 12099 13574 12111 13626
rect 12163 13574 12175 13626
rect 12227 13574 12239 13626
rect 12291 13574 12303 13626
rect 12355 13574 16486 13626
rect 16538 13574 16550 13626
rect 16602 13574 16614 13626
rect 16666 13574 16678 13626
rect 16730 13574 16742 13626
rect 16794 13574 18860 13626
rect 1104 13552 18860 13574
rect 1104 13082 19019 13104
rect 1104 13030 5388 13082
rect 5440 13030 5452 13082
rect 5504 13030 5516 13082
rect 5568 13030 5580 13082
rect 5632 13030 5644 13082
rect 5696 13030 9827 13082
rect 9879 13030 9891 13082
rect 9943 13030 9955 13082
rect 10007 13030 10019 13082
rect 10071 13030 10083 13082
rect 10135 13030 14266 13082
rect 14318 13030 14330 13082
rect 14382 13030 14394 13082
rect 14446 13030 14458 13082
rect 14510 13030 14522 13082
rect 14574 13030 18705 13082
rect 18757 13030 18769 13082
rect 18821 13030 18833 13082
rect 18885 13030 18897 13082
rect 18949 13030 18961 13082
rect 19013 13030 19019 13082
rect 1104 13008 19019 13030
rect 1104 12538 18860 12560
rect 1104 12486 3169 12538
rect 3221 12486 3233 12538
rect 3285 12486 3297 12538
rect 3349 12486 3361 12538
rect 3413 12486 3425 12538
rect 3477 12486 7608 12538
rect 7660 12486 7672 12538
rect 7724 12486 7736 12538
rect 7788 12486 7800 12538
rect 7852 12486 7864 12538
rect 7916 12486 12047 12538
rect 12099 12486 12111 12538
rect 12163 12486 12175 12538
rect 12227 12486 12239 12538
rect 12291 12486 12303 12538
rect 12355 12486 16486 12538
rect 16538 12486 16550 12538
rect 16602 12486 16614 12538
rect 16666 12486 16678 12538
rect 16730 12486 16742 12538
rect 16794 12486 18860 12538
rect 1104 12464 18860 12486
rect 1104 11994 19019 12016
rect 1104 11942 5388 11994
rect 5440 11942 5452 11994
rect 5504 11942 5516 11994
rect 5568 11942 5580 11994
rect 5632 11942 5644 11994
rect 5696 11942 9827 11994
rect 9879 11942 9891 11994
rect 9943 11942 9955 11994
rect 10007 11942 10019 11994
rect 10071 11942 10083 11994
rect 10135 11942 14266 11994
rect 14318 11942 14330 11994
rect 14382 11942 14394 11994
rect 14446 11942 14458 11994
rect 14510 11942 14522 11994
rect 14574 11942 18705 11994
rect 18757 11942 18769 11994
rect 18821 11942 18833 11994
rect 18885 11942 18897 11994
rect 18949 11942 18961 11994
rect 19013 11942 19019 11994
rect 1104 11920 19019 11942
rect 1104 11450 18860 11472
rect 1104 11398 3169 11450
rect 3221 11398 3233 11450
rect 3285 11398 3297 11450
rect 3349 11398 3361 11450
rect 3413 11398 3425 11450
rect 3477 11398 7608 11450
rect 7660 11398 7672 11450
rect 7724 11398 7736 11450
rect 7788 11398 7800 11450
rect 7852 11398 7864 11450
rect 7916 11398 12047 11450
rect 12099 11398 12111 11450
rect 12163 11398 12175 11450
rect 12227 11398 12239 11450
rect 12291 11398 12303 11450
rect 12355 11398 16486 11450
rect 16538 11398 16550 11450
rect 16602 11398 16614 11450
rect 16666 11398 16678 11450
rect 16730 11398 16742 11450
rect 16794 11398 18860 11450
rect 1104 11376 18860 11398
rect 1104 10906 19019 10928
rect 1104 10854 5388 10906
rect 5440 10854 5452 10906
rect 5504 10854 5516 10906
rect 5568 10854 5580 10906
rect 5632 10854 5644 10906
rect 5696 10854 9827 10906
rect 9879 10854 9891 10906
rect 9943 10854 9955 10906
rect 10007 10854 10019 10906
rect 10071 10854 10083 10906
rect 10135 10854 14266 10906
rect 14318 10854 14330 10906
rect 14382 10854 14394 10906
rect 14446 10854 14458 10906
rect 14510 10854 14522 10906
rect 14574 10854 18705 10906
rect 18757 10854 18769 10906
rect 18821 10854 18833 10906
rect 18885 10854 18897 10906
rect 18949 10854 18961 10906
rect 19013 10854 19019 10906
rect 1104 10832 19019 10854
rect 1104 10362 18860 10384
rect 1104 10310 3169 10362
rect 3221 10310 3233 10362
rect 3285 10310 3297 10362
rect 3349 10310 3361 10362
rect 3413 10310 3425 10362
rect 3477 10310 7608 10362
rect 7660 10310 7672 10362
rect 7724 10310 7736 10362
rect 7788 10310 7800 10362
rect 7852 10310 7864 10362
rect 7916 10310 12047 10362
rect 12099 10310 12111 10362
rect 12163 10310 12175 10362
rect 12227 10310 12239 10362
rect 12291 10310 12303 10362
rect 12355 10310 16486 10362
rect 16538 10310 16550 10362
rect 16602 10310 16614 10362
rect 16666 10310 16678 10362
rect 16730 10310 16742 10362
rect 16794 10310 18860 10362
rect 1104 10288 18860 10310
rect 1104 9818 19019 9840
rect 1104 9766 5388 9818
rect 5440 9766 5452 9818
rect 5504 9766 5516 9818
rect 5568 9766 5580 9818
rect 5632 9766 5644 9818
rect 5696 9766 9827 9818
rect 9879 9766 9891 9818
rect 9943 9766 9955 9818
rect 10007 9766 10019 9818
rect 10071 9766 10083 9818
rect 10135 9766 14266 9818
rect 14318 9766 14330 9818
rect 14382 9766 14394 9818
rect 14446 9766 14458 9818
rect 14510 9766 14522 9818
rect 14574 9766 18705 9818
rect 18757 9766 18769 9818
rect 18821 9766 18833 9818
rect 18885 9766 18897 9818
rect 18949 9766 18961 9818
rect 19013 9766 19019 9818
rect 1104 9744 19019 9766
rect 18506 9324 18512 9376
rect 18564 9324 18570 9376
rect 1104 9274 18860 9296
rect 1104 9222 3169 9274
rect 3221 9222 3233 9274
rect 3285 9222 3297 9274
rect 3349 9222 3361 9274
rect 3413 9222 3425 9274
rect 3477 9222 7608 9274
rect 7660 9222 7672 9274
rect 7724 9222 7736 9274
rect 7788 9222 7800 9274
rect 7852 9222 7864 9274
rect 7916 9222 12047 9274
rect 12099 9222 12111 9274
rect 12163 9222 12175 9274
rect 12227 9222 12239 9274
rect 12291 9222 12303 9274
rect 12355 9222 16486 9274
rect 16538 9222 16550 9274
rect 16602 9222 16614 9274
rect 16666 9222 16678 9274
rect 16730 9222 16742 9274
rect 16794 9222 18860 9274
rect 1104 9200 18860 9222
rect 1104 8730 19019 8752
rect 1104 8678 5388 8730
rect 5440 8678 5452 8730
rect 5504 8678 5516 8730
rect 5568 8678 5580 8730
rect 5632 8678 5644 8730
rect 5696 8678 9827 8730
rect 9879 8678 9891 8730
rect 9943 8678 9955 8730
rect 10007 8678 10019 8730
rect 10071 8678 10083 8730
rect 10135 8678 14266 8730
rect 14318 8678 14330 8730
rect 14382 8678 14394 8730
rect 14446 8678 14458 8730
rect 14510 8678 14522 8730
rect 14574 8678 18705 8730
rect 18757 8678 18769 8730
rect 18821 8678 18833 8730
rect 18885 8678 18897 8730
rect 18949 8678 18961 8730
rect 19013 8678 19019 8730
rect 1104 8656 19019 8678
rect 18414 8576 18420 8628
rect 18472 8576 18478 8628
rect 15933 8551 15991 8557
rect 15933 8517 15945 8551
rect 15979 8548 15991 8551
rect 16942 8548 16948 8560
rect 15979 8520 16948 8548
rect 15979 8517 15991 8520
rect 15933 8511 15991 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 16025 8483 16083 8489
rect 16025 8449 16037 8483
rect 16071 8480 16083 8483
rect 17126 8480 17132 8492
rect 16071 8452 17132 8480
rect 16071 8449 16083 8452
rect 16025 8443 16083 8449
rect 15764 8412 15792 8443
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 15930 8412 15936 8424
rect 15764 8384 15936 8412
rect 15930 8372 15936 8384
rect 15988 8372 15994 8424
rect 15746 8304 15752 8356
rect 15804 8304 15810 8356
rect 1104 8186 18860 8208
rect 1104 8134 3169 8186
rect 3221 8134 3233 8186
rect 3285 8134 3297 8186
rect 3349 8134 3361 8186
rect 3413 8134 3425 8186
rect 3477 8134 7608 8186
rect 7660 8134 7672 8186
rect 7724 8134 7736 8186
rect 7788 8134 7800 8186
rect 7852 8134 7864 8186
rect 7916 8134 12047 8186
rect 12099 8134 12111 8186
rect 12163 8134 12175 8186
rect 12227 8134 12239 8186
rect 12291 8134 12303 8186
rect 12355 8134 16486 8186
rect 16538 8134 16550 8186
rect 16602 8134 16614 8186
rect 16666 8134 16678 8186
rect 16730 8134 16742 8186
rect 16794 8134 18860 8186
rect 1104 8112 18860 8134
rect 17034 8072 17040 8084
rect 15856 8044 17040 8072
rect 15856 7877 15884 8044
rect 17034 8032 17040 8044
rect 17092 8032 17098 8084
rect 15930 7964 15936 8016
rect 15988 8004 15994 8016
rect 16025 8007 16083 8013
rect 16025 8004 16037 8007
rect 15988 7976 16037 8004
rect 15988 7964 15994 7976
rect 16025 7973 16037 7976
rect 16071 8004 16083 8007
rect 16390 8004 16396 8016
rect 16071 7976 16396 8004
rect 16071 7973 16083 7976
rect 16025 7967 16083 7973
rect 16390 7964 16396 7976
rect 16448 8004 16454 8016
rect 16448 7976 17724 8004
rect 16448 7964 16454 7976
rect 16942 7896 16948 7948
rect 17000 7936 17006 7948
rect 17405 7939 17463 7945
rect 17405 7936 17417 7939
rect 17000 7908 17417 7936
rect 17000 7896 17006 7908
rect 17405 7905 17417 7908
rect 17451 7905 17463 7939
rect 17405 7899 17463 7905
rect 15841 7871 15899 7877
rect 15841 7868 15853 7871
rect 15672 7840 15853 7868
rect 14918 7692 14924 7744
rect 14976 7732 14982 7744
rect 15672 7741 15700 7840
rect 15841 7837 15853 7840
rect 15887 7837 15899 7871
rect 15841 7831 15899 7837
rect 16758 7828 16764 7880
rect 16816 7828 16822 7880
rect 17696 7877 17724 7976
rect 18414 7896 18420 7948
rect 18472 7896 18478 7948
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17773 7871 17831 7877
rect 17773 7837 17785 7871
rect 17819 7868 17831 7871
rect 17819 7840 17908 7868
rect 17819 7837 17831 7840
rect 17773 7831 17831 7837
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 14976 7704 15669 7732
rect 14976 7692 14982 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 16114 7692 16120 7744
rect 16172 7692 16178 7744
rect 17402 7692 17408 7744
rect 17460 7692 17466 7744
rect 17586 7692 17592 7744
rect 17644 7692 17650 7744
rect 17880 7741 17908 7840
rect 17865 7735 17923 7741
rect 17865 7701 17877 7735
rect 17911 7732 17923 7735
rect 18138 7732 18144 7744
rect 17911 7704 18144 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18138 7692 18144 7704
rect 18196 7692 18202 7744
rect 1104 7642 19019 7664
rect 1104 7590 5388 7642
rect 5440 7590 5452 7642
rect 5504 7590 5516 7642
rect 5568 7590 5580 7642
rect 5632 7590 5644 7642
rect 5696 7590 9827 7642
rect 9879 7590 9891 7642
rect 9943 7590 9955 7642
rect 10007 7590 10019 7642
rect 10071 7590 10083 7642
rect 10135 7590 14266 7642
rect 14318 7590 14330 7642
rect 14382 7590 14394 7642
rect 14446 7590 14458 7642
rect 14510 7590 14522 7642
rect 14574 7590 18705 7642
rect 18757 7590 18769 7642
rect 18821 7590 18833 7642
rect 18885 7590 18897 7642
rect 18949 7590 18961 7642
rect 19013 7590 19019 7642
rect 1104 7568 19019 7590
rect 14918 7488 14924 7540
rect 14976 7488 14982 7540
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18414 7528 18420 7540
rect 18371 7500 18420 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 16045 7395 16103 7401
rect 16045 7361 16057 7395
rect 16091 7392 16103 7395
rect 16132 7392 16160 7488
rect 16945 7395 17003 7401
rect 16945 7392 16957 7395
rect 16091 7364 16160 7392
rect 16546 7364 16957 7392
rect 16091 7361 16103 7364
rect 16045 7355 16103 7361
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16546 7324 16574 7364
rect 16945 7361 16957 7364
rect 16991 7361 17003 7395
rect 16945 7355 17003 7361
rect 17212 7395 17270 7401
rect 17212 7361 17224 7395
rect 17258 7392 17270 7395
rect 17586 7392 17592 7404
rect 17258 7364 17592 7392
rect 17258 7361 17270 7364
rect 17212 7355 17270 7361
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 16347 7296 16574 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16114 7148 16120 7200
rect 16172 7188 16178 7200
rect 16316 7188 16344 7287
rect 16172 7160 16344 7188
rect 16172 7148 16178 7160
rect 1104 7098 18860 7120
rect 1104 7046 3169 7098
rect 3221 7046 3233 7098
rect 3285 7046 3297 7098
rect 3349 7046 3361 7098
rect 3413 7046 3425 7098
rect 3477 7046 7608 7098
rect 7660 7046 7672 7098
rect 7724 7046 7736 7098
rect 7788 7046 7800 7098
rect 7852 7046 7864 7098
rect 7916 7046 12047 7098
rect 12099 7046 12111 7098
rect 12163 7046 12175 7098
rect 12227 7046 12239 7098
rect 12291 7046 12303 7098
rect 12355 7046 16486 7098
rect 16538 7046 16550 7098
rect 16602 7046 16614 7098
rect 16666 7046 16678 7098
rect 16730 7046 16742 7098
rect 16794 7046 18860 7098
rect 1104 7024 18860 7046
rect 16390 6944 16396 6996
rect 16448 6944 16454 6996
rect 16592 6956 17080 6984
rect 16408 6916 16436 6944
rect 16592 6916 16620 6956
rect 16942 6916 16948 6928
rect 16408 6888 16620 6916
rect 15657 6851 15715 6857
rect 15657 6848 15669 6851
rect 15396 6820 15669 6848
rect 15396 6789 15424 6820
rect 15657 6817 15669 6820
rect 15703 6817 15715 6851
rect 15657 6811 15715 6817
rect 15746 6808 15752 6860
rect 15804 6848 15810 6860
rect 16592 6857 16620 6888
rect 16776 6888 16948 6916
rect 16776 6857 16804 6888
rect 16942 6876 16948 6888
rect 17000 6876 17006 6928
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 15804 6820 16221 6848
rect 15804 6808 15810 6820
rect 16209 6817 16221 6820
rect 16255 6817 16267 6851
rect 16209 6811 16267 6817
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 16577 6851 16635 6857
rect 16577 6817 16589 6851
rect 16623 6817 16635 6851
rect 16577 6811 16635 6817
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6848 16819 6851
rect 17052 6848 17080 6956
rect 17402 6944 17408 6996
rect 17460 6944 17466 6996
rect 17586 6944 17592 6996
rect 17644 6944 17650 6996
rect 17678 6876 17684 6928
rect 17736 6916 17742 6928
rect 17736 6888 18000 6916
rect 17736 6876 17742 6888
rect 17972 6857 18000 6888
rect 17865 6851 17923 6857
rect 17865 6848 17877 6851
rect 16807 6820 16841 6848
rect 17052 6820 17877 6848
rect 16807 6817 16819 6820
rect 16761 6811 16819 6817
rect 17865 6817 17877 6820
rect 17911 6817 17923 6851
rect 17865 6811 17923 6817
rect 17957 6851 18015 6857
rect 17957 6817 17969 6851
rect 18003 6848 18015 6851
rect 18003 6820 18037 6848
rect 18003 6817 18015 6820
rect 17957 6811 18015 6817
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 15565 6783 15623 6789
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 16408 6780 16436 6811
rect 18138 6808 18144 6860
rect 18196 6808 18202 6860
rect 15611 6752 16436 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 16666 6740 16672 6792
rect 16724 6740 16730 6792
rect 16853 6783 16911 6789
rect 16853 6749 16865 6783
rect 16899 6780 16911 6783
rect 17037 6783 17095 6789
rect 17037 6780 17049 6783
rect 16899 6752 17049 6780
rect 16899 6749 16911 6752
rect 16853 6743 16911 6749
rect 17037 6749 17049 6752
rect 17083 6749 17095 6783
rect 17037 6743 17095 6749
rect 16022 6672 16028 6724
rect 16080 6712 16086 6724
rect 16868 6712 16896 6743
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 18049 6783 18107 6789
rect 18049 6780 18061 6783
rect 17184 6752 18061 6780
rect 17184 6740 17190 6752
rect 18049 6749 18061 6752
rect 18095 6749 18107 6783
rect 18049 6743 18107 6749
rect 16080 6684 16896 6712
rect 16080 6672 16086 6684
rect 15473 6647 15531 6653
rect 15473 6613 15485 6647
rect 15519 6644 15531 6647
rect 16850 6644 16856 6656
rect 15519 6616 16856 6644
rect 15519 6613 15531 6616
rect 15473 6607 15531 6613
rect 16850 6604 16856 6616
rect 16908 6604 16914 6656
rect 17405 6647 17463 6653
rect 17405 6613 17417 6647
rect 17451 6644 17463 6647
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17451 6616 17693 6644
rect 17451 6613 17463 6616
rect 17405 6607 17463 6613
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 1104 6554 19019 6576
rect 1104 6502 5388 6554
rect 5440 6502 5452 6554
rect 5504 6502 5516 6554
rect 5568 6502 5580 6554
rect 5632 6502 5644 6554
rect 5696 6502 9827 6554
rect 9879 6502 9891 6554
rect 9943 6502 9955 6554
rect 10007 6502 10019 6554
rect 10071 6502 10083 6554
rect 10135 6502 14266 6554
rect 14318 6502 14330 6554
rect 14382 6502 14394 6554
rect 14446 6502 14458 6554
rect 14510 6502 14522 6554
rect 14574 6502 18705 6554
rect 18757 6502 18769 6554
rect 18821 6502 18833 6554
rect 18885 6502 18897 6554
rect 18949 6502 18961 6554
rect 19013 6502 19019 6554
rect 1104 6480 19019 6502
rect 16666 6400 16672 6452
rect 16724 6440 16730 6452
rect 17218 6440 17224 6452
rect 16724 6412 17224 6440
rect 16724 6400 16730 6412
rect 17218 6400 17224 6412
rect 17276 6400 17282 6452
rect 1104 6010 18860 6032
rect 1104 5958 3169 6010
rect 3221 5958 3233 6010
rect 3285 5958 3297 6010
rect 3349 5958 3361 6010
rect 3413 5958 3425 6010
rect 3477 5958 7608 6010
rect 7660 5958 7672 6010
rect 7724 5958 7736 6010
rect 7788 5958 7800 6010
rect 7852 5958 7864 6010
rect 7916 5958 12047 6010
rect 12099 5958 12111 6010
rect 12163 5958 12175 6010
rect 12227 5958 12239 6010
rect 12291 5958 12303 6010
rect 12355 5958 16486 6010
rect 16538 5958 16550 6010
rect 16602 5958 16614 6010
rect 16666 5958 16678 6010
rect 16730 5958 16742 6010
rect 16794 5958 18860 6010
rect 1104 5936 18860 5958
rect 16114 5856 16120 5908
rect 16172 5856 16178 5908
rect 17402 5584 17408 5636
rect 17460 5584 17466 5636
rect 1104 5466 19019 5488
rect 1104 5414 5388 5466
rect 5440 5414 5452 5466
rect 5504 5414 5516 5466
rect 5568 5414 5580 5466
rect 5632 5414 5644 5466
rect 5696 5414 9827 5466
rect 9879 5414 9891 5466
rect 9943 5414 9955 5466
rect 10007 5414 10019 5466
rect 10071 5414 10083 5466
rect 10135 5414 14266 5466
rect 14318 5414 14330 5466
rect 14382 5414 14394 5466
rect 14446 5414 14458 5466
rect 14510 5414 14522 5466
rect 14574 5414 18705 5466
rect 18757 5414 18769 5466
rect 18821 5414 18833 5466
rect 18885 5414 18897 5466
rect 18949 5414 18961 5466
rect 19013 5414 19019 5466
rect 1104 5392 19019 5414
rect 16117 5355 16175 5361
rect 16117 5321 16129 5355
rect 16163 5352 16175 5355
rect 16390 5352 16396 5364
rect 16163 5324 16396 5352
rect 16163 5321 16175 5324
rect 16117 5315 16175 5321
rect 16390 5312 16396 5324
rect 16448 5352 16454 5364
rect 17034 5352 17040 5364
rect 16448 5324 17040 5352
rect 16448 5312 16454 5324
rect 17034 5312 17040 5324
rect 17092 5312 17098 5364
rect 15933 5287 15991 5293
rect 15933 5253 15945 5287
rect 15979 5284 15991 5287
rect 16022 5284 16028 5296
rect 15979 5256 16028 5284
rect 15979 5253 15991 5256
rect 15933 5247 15991 5253
rect 16022 5244 16028 5256
rect 16080 5244 16086 5296
rect 16209 5219 16267 5225
rect 16209 5185 16221 5219
rect 16255 5216 16267 5219
rect 16298 5216 16304 5228
rect 16255 5188 16304 5216
rect 16255 5185 16267 5188
rect 16209 5179 16267 5185
rect 16298 5176 16304 5188
rect 16356 5216 16362 5228
rect 16669 5219 16727 5225
rect 16356 5188 16574 5216
rect 16356 5176 16362 5188
rect 16546 5148 16574 5188
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16850 5216 16856 5228
rect 16715 5188 16856 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 17678 5148 17684 5160
rect 16546 5120 17684 5148
rect 17678 5108 17684 5120
rect 17736 5108 17742 5160
rect 15930 4972 15936 5024
rect 15988 4972 15994 5024
rect 17402 4972 17408 5024
rect 17460 5012 17466 5024
rect 17957 5015 18015 5021
rect 17957 5012 17969 5015
rect 17460 4984 17969 5012
rect 17460 4972 17466 4984
rect 17957 4981 17969 4984
rect 18003 4981 18015 5015
rect 17957 4975 18015 4981
rect 1104 4922 18860 4944
rect 1104 4870 3169 4922
rect 3221 4870 3233 4922
rect 3285 4870 3297 4922
rect 3349 4870 3361 4922
rect 3413 4870 3425 4922
rect 3477 4870 7608 4922
rect 7660 4870 7672 4922
rect 7724 4870 7736 4922
rect 7788 4870 7800 4922
rect 7852 4870 7864 4922
rect 7916 4870 12047 4922
rect 12099 4870 12111 4922
rect 12163 4870 12175 4922
rect 12227 4870 12239 4922
rect 12291 4870 12303 4922
rect 12355 4870 16486 4922
rect 16538 4870 16550 4922
rect 16602 4870 16614 4922
rect 16666 4870 16678 4922
rect 16730 4870 16742 4922
rect 16794 4870 18860 4922
rect 1104 4848 18860 4870
rect 15749 4607 15807 4613
rect 15749 4573 15761 4607
rect 15795 4604 15807 4607
rect 15795 4576 16160 4604
rect 15795 4573 15807 4576
rect 15749 4567 15807 4573
rect 16022 4545 16028 4548
rect 16016 4499 16028 4545
rect 16022 4496 16028 4499
rect 16080 4496 16086 4548
rect 16132 4480 16160 4576
rect 17310 4564 17316 4616
rect 17368 4564 17374 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17678 4604 17684 4616
rect 17635 4576 17684 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 17678 4564 17684 4576
rect 17736 4564 17742 4616
rect 16114 4428 16120 4480
rect 16172 4428 16178 4480
rect 17126 4428 17132 4480
rect 17184 4428 17190 4480
rect 1104 4378 19019 4400
rect 1104 4326 5388 4378
rect 5440 4326 5452 4378
rect 5504 4326 5516 4378
rect 5568 4326 5580 4378
rect 5632 4326 5644 4378
rect 5696 4326 9827 4378
rect 9879 4326 9891 4378
rect 9943 4326 9955 4378
rect 10007 4326 10019 4378
rect 10071 4326 10083 4378
rect 10135 4326 14266 4378
rect 14318 4326 14330 4378
rect 14382 4326 14394 4378
rect 14446 4326 14458 4378
rect 14510 4326 14522 4378
rect 14574 4326 18705 4378
rect 18757 4326 18769 4378
rect 18821 4326 18833 4378
rect 18885 4326 18897 4378
rect 18949 4326 18961 4378
rect 19013 4326 19019 4378
rect 1104 4304 19019 4326
rect 15933 4267 15991 4273
rect 15933 4233 15945 4267
rect 15979 4264 15991 4267
rect 16022 4264 16028 4276
rect 15979 4236 16028 4264
rect 15979 4233 15991 4236
rect 15933 4227 15991 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 15930 4088 15936 4140
rect 15988 4128 15994 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15988 4100 16129 4128
rect 15988 4088 15994 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 16117 4091 16175 4097
rect 16298 4088 16304 4140
rect 16356 4088 16362 4140
rect 16390 4088 16396 4140
rect 16448 4088 16454 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17678 4128 17684 4140
rect 17359 4100 17684 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17678 4088 17684 4100
rect 17736 4088 17742 4140
rect 18322 4020 18328 4072
rect 18380 4020 18386 4072
rect 1104 3834 18860 3856
rect 1104 3782 3169 3834
rect 3221 3782 3233 3834
rect 3285 3782 3297 3834
rect 3349 3782 3361 3834
rect 3413 3782 3425 3834
rect 3477 3782 7608 3834
rect 7660 3782 7672 3834
rect 7724 3782 7736 3834
rect 7788 3782 7800 3834
rect 7852 3782 7864 3834
rect 7916 3782 12047 3834
rect 12099 3782 12111 3834
rect 12163 3782 12175 3834
rect 12227 3782 12239 3834
rect 12291 3782 12303 3834
rect 12355 3782 16486 3834
rect 16538 3782 16550 3834
rect 16602 3782 16614 3834
rect 16666 3782 16678 3834
rect 16730 3782 16742 3834
rect 16794 3782 18860 3834
rect 1104 3760 18860 3782
rect 17310 3680 17316 3732
rect 17368 3720 17374 3732
rect 17497 3723 17555 3729
rect 17497 3720 17509 3723
rect 17368 3692 17509 3720
rect 17368 3680 17374 3692
rect 17497 3689 17509 3692
rect 17543 3689 17555 3723
rect 17497 3683 17555 3689
rect 16390 3612 16396 3664
rect 16448 3652 16454 3664
rect 18233 3655 18291 3661
rect 18233 3652 18245 3655
rect 16448 3624 18245 3652
rect 16448 3612 16454 3624
rect 18233 3621 18245 3624
rect 18279 3621 18291 3655
rect 18233 3615 18291 3621
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 18049 3587 18107 3593
rect 18049 3584 18061 3587
rect 17184 3556 18061 3584
rect 17184 3544 17190 3556
rect 18049 3553 18061 3556
rect 18095 3553 18107 3587
rect 18049 3547 18107 3553
rect 4982 3476 4988 3528
rect 5040 3516 5046 3528
rect 16850 3516 16856 3528
rect 5040 3488 16856 3516
rect 5040 3476 5046 3488
rect 16850 3476 16856 3488
rect 16908 3476 16914 3528
rect 17402 3476 17408 3528
rect 17460 3476 17466 3528
rect 18414 3408 18420 3460
rect 18472 3408 18478 3460
rect 16114 3340 16120 3392
rect 16172 3380 16178 3392
rect 16482 3380 16488 3392
rect 16172 3352 16488 3380
rect 16172 3340 16178 3352
rect 16482 3340 16488 3352
rect 16540 3340 16546 3392
rect 1104 3290 19019 3312
rect 1104 3238 5388 3290
rect 5440 3238 5452 3290
rect 5504 3238 5516 3290
rect 5568 3238 5580 3290
rect 5632 3238 5644 3290
rect 5696 3238 9827 3290
rect 9879 3238 9891 3290
rect 9943 3238 9955 3290
rect 10007 3238 10019 3290
rect 10071 3238 10083 3290
rect 10135 3238 14266 3290
rect 14318 3238 14330 3290
rect 14382 3238 14394 3290
rect 14446 3238 14458 3290
rect 14510 3238 14522 3290
rect 14574 3238 18705 3290
rect 18757 3238 18769 3290
rect 18821 3238 18833 3290
rect 18885 3238 18897 3290
rect 18949 3238 18961 3290
rect 19013 3238 19019 3290
rect 1104 3216 19019 3238
rect 16408 3148 16574 3176
rect 16408 3117 16436 3148
rect 16393 3111 16451 3117
rect 16393 3077 16405 3111
rect 16439 3077 16451 3111
rect 16546 3108 16574 3148
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 17736 3148 18061 3176
rect 17736 3136 17742 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 16914 3111 16972 3117
rect 16914 3108 16926 3111
rect 16546 3080 16926 3108
rect 16393 3071 16451 3077
rect 16914 3077 16926 3080
rect 16960 3077 16972 3111
rect 16914 3071 16972 3077
rect 16206 3000 16212 3052
rect 16264 3000 16270 3052
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16485 3043 16543 3049
rect 16485 3040 16497 3043
rect 16408 3012 16497 3040
rect 16224 2972 16252 3000
rect 16408 2972 16436 3012
rect 16485 3009 16497 3012
rect 16531 3009 16543 3043
rect 16485 3003 16543 3009
rect 16669 2975 16727 2981
rect 16669 2972 16681 2975
rect 16224 2944 16436 2972
rect 16546 2944 16681 2972
rect 16546 2916 16574 2944
rect 16669 2941 16681 2944
rect 16715 2941 16727 2975
rect 16669 2935 16727 2941
rect 16482 2864 16488 2916
rect 16540 2876 16574 2916
rect 16540 2864 16546 2876
rect 1104 2746 18860 2768
rect 1104 2694 3169 2746
rect 3221 2694 3233 2746
rect 3285 2694 3297 2746
rect 3349 2694 3361 2746
rect 3413 2694 3425 2746
rect 3477 2694 7608 2746
rect 7660 2694 7672 2746
rect 7724 2694 7736 2746
rect 7788 2694 7800 2746
rect 7852 2694 7864 2746
rect 7916 2694 12047 2746
rect 12099 2694 12111 2746
rect 12163 2694 12175 2746
rect 12227 2694 12239 2746
rect 12291 2694 12303 2746
rect 12355 2694 16486 2746
rect 16538 2694 16550 2746
rect 16602 2694 16614 2746
rect 16666 2694 16678 2746
rect 16730 2694 16742 2746
rect 16794 2694 18860 2746
rect 1104 2672 18860 2694
rect 15197 2635 15255 2641
rect 15197 2601 15209 2635
rect 15243 2632 15255 2635
rect 16206 2632 16212 2644
rect 15243 2604 16212 2632
rect 15243 2601 15255 2604
rect 15197 2595 15255 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 18509 2635 18567 2641
rect 18509 2632 18521 2635
rect 18472 2604 18521 2632
rect 18472 2592 18478 2604
rect 18509 2601 18521 2604
rect 18555 2601 18567 2635
rect 18509 2595 18567 2601
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17865 2499 17923 2505
rect 17865 2496 17877 2499
rect 17736 2468 17877 2496
rect 17736 2456 17742 2468
rect 17865 2465 17877 2468
rect 17911 2465 17923 2499
rect 17865 2459 17923 2465
rect 15010 2388 15016 2440
rect 15068 2388 15074 2440
rect 1104 2202 19019 2224
rect 1104 2150 5388 2202
rect 5440 2150 5452 2202
rect 5504 2150 5516 2202
rect 5568 2150 5580 2202
rect 5632 2150 5644 2202
rect 5696 2150 9827 2202
rect 9879 2150 9891 2202
rect 9943 2150 9955 2202
rect 10007 2150 10019 2202
rect 10071 2150 10083 2202
rect 10135 2150 14266 2202
rect 14318 2150 14330 2202
rect 14382 2150 14394 2202
rect 14446 2150 14458 2202
rect 14510 2150 14522 2202
rect 14574 2150 18705 2202
rect 18757 2150 18769 2202
rect 18821 2150 18833 2202
rect 18885 2150 18897 2202
rect 18949 2150 18961 2202
rect 19013 2150 19019 2202
rect 1104 2128 19019 2150
<< via1 >>
rect 3169 47302 3221 47354
rect 3233 47302 3285 47354
rect 3297 47302 3349 47354
rect 3361 47302 3413 47354
rect 3425 47302 3477 47354
rect 7608 47302 7660 47354
rect 7672 47302 7724 47354
rect 7736 47302 7788 47354
rect 7800 47302 7852 47354
rect 7864 47302 7916 47354
rect 12047 47302 12099 47354
rect 12111 47302 12163 47354
rect 12175 47302 12227 47354
rect 12239 47302 12291 47354
rect 12303 47302 12355 47354
rect 16486 47302 16538 47354
rect 16550 47302 16602 47354
rect 16614 47302 16666 47354
rect 16678 47302 16730 47354
rect 16742 47302 16794 47354
rect 18512 47243 18564 47252
rect 18512 47209 18521 47243
rect 18521 47209 18555 47243
rect 18555 47209 18564 47243
rect 18512 47200 18564 47209
rect 5388 46758 5440 46810
rect 5452 46758 5504 46810
rect 5516 46758 5568 46810
rect 5580 46758 5632 46810
rect 5644 46758 5696 46810
rect 9827 46758 9879 46810
rect 9891 46758 9943 46810
rect 9955 46758 10007 46810
rect 10019 46758 10071 46810
rect 10083 46758 10135 46810
rect 14266 46758 14318 46810
rect 14330 46758 14382 46810
rect 14394 46758 14446 46810
rect 14458 46758 14510 46810
rect 14522 46758 14574 46810
rect 18705 46758 18757 46810
rect 18769 46758 18821 46810
rect 18833 46758 18885 46810
rect 18897 46758 18949 46810
rect 18961 46758 19013 46810
rect 3169 46214 3221 46266
rect 3233 46214 3285 46266
rect 3297 46214 3349 46266
rect 3361 46214 3413 46266
rect 3425 46214 3477 46266
rect 7608 46214 7660 46266
rect 7672 46214 7724 46266
rect 7736 46214 7788 46266
rect 7800 46214 7852 46266
rect 7864 46214 7916 46266
rect 12047 46214 12099 46266
rect 12111 46214 12163 46266
rect 12175 46214 12227 46266
rect 12239 46214 12291 46266
rect 12303 46214 12355 46266
rect 16486 46214 16538 46266
rect 16550 46214 16602 46266
rect 16614 46214 16666 46266
rect 16678 46214 16730 46266
rect 16742 46214 16794 46266
rect 5388 45670 5440 45722
rect 5452 45670 5504 45722
rect 5516 45670 5568 45722
rect 5580 45670 5632 45722
rect 5644 45670 5696 45722
rect 9827 45670 9879 45722
rect 9891 45670 9943 45722
rect 9955 45670 10007 45722
rect 10019 45670 10071 45722
rect 10083 45670 10135 45722
rect 14266 45670 14318 45722
rect 14330 45670 14382 45722
rect 14394 45670 14446 45722
rect 14458 45670 14510 45722
rect 14522 45670 14574 45722
rect 18705 45670 18757 45722
rect 18769 45670 18821 45722
rect 18833 45670 18885 45722
rect 18897 45670 18949 45722
rect 18961 45670 19013 45722
rect 3169 45126 3221 45178
rect 3233 45126 3285 45178
rect 3297 45126 3349 45178
rect 3361 45126 3413 45178
rect 3425 45126 3477 45178
rect 7608 45126 7660 45178
rect 7672 45126 7724 45178
rect 7736 45126 7788 45178
rect 7800 45126 7852 45178
rect 7864 45126 7916 45178
rect 12047 45126 12099 45178
rect 12111 45126 12163 45178
rect 12175 45126 12227 45178
rect 12239 45126 12291 45178
rect 12303 45126 12355 45178
rect 16486 45126 16538 45178
rect 16550 45126 16602 45178
rect 16614 45126 16666 45178
rect 16678 45126 16730 45178
rect 16742 45126 16794 45178
rect 5388 44582 5440 44634
rect 5452 44582 5504 44634
rect 5516 44582 5568 44634
rect 5580 44582 5632 44634
rect 5644 44582 5696 44634
rect 9827 44582 9879 44634
rect 9891 44582 9943 44634
rect 9955 44582 10007 44634
rect 10019 44582 10071 44634
rect 10083 44582 10135 44634
rect 14266 44582 14318 44634
rect 14330 44582 14382 44634
rect 14394 44582 14446 44634
rect 14458 44582 14510 44634
rect 14522 44582 14574 44634
rect 18705 44582 18757 44634
rect 18769 44582 18821 44634
rect 18833 44582 18885 44634
rect 18897 44582 18949 44634
rect 18961 44582 19013 44634
rect 3169 44038 3221 44090
rect 3233 44038 3285 44090
rect 3297 44038 3349 44090
rect 3361 44038 3413 44090
rect 3425 44038 3477 44090
rect 7608 44038 7660 44090
rect 7672 44038 7724 44090
rect 7736 44038 7788 44090
rect 7800 44038 7852 44090
rect 7864 44038 7916 44090
rect 12047 44038 12099 44090
rect 12111 44038 12163 44090
rect 12175 44038 12227 44090
rect 12239 44038 12291 44090
rect 12303 44038 12355 44090
rect 16486 44038 16538 44090
rect 16550 44038 16602 44090
rect 16614 44038 16666 44090
rect 16678 44038 16730 44090
rect 16742 44038 16794 44090
rect 5388 43494 5440 43546
rect 5452 43494 5504 43546
rect 5516 43494 5568 43546
rect 5580 43494 5632 43546
rect 5644 43494 5696 43546
rect 9827 43494 9879 43546
rect 9891 43494 9943 43546
rect 9955 43494 10007 43546
rect 10019 43494 10071 43546
rect 10083 43494 10135 43546
rect 14266 43494 14318 43546
rect 14330 43494 14382 43546
rect 14394 43494 14446 43546
rect 14458 43494 14510 43546
rect 14522 43494 14574 43546
rect 18705 43494 18757 43546
rect 18769 43494 18821 43546
rect 18833 43494 18885 43546
rect 18897 43494 18949 43546
rect 18961 43494 19013 43546
rect 3169 42950 3221 43002
rect 3233 42950 3285 43002
rect 3297 42950 3349 43002
rect 3361 42950 3413 43002
rect 3425 42950 3477 43002
rect 7608 42950 7660 43002
rect 7672 42950 7724 43002
rect 7736 42950 7788 43002
rect 7800 42950 7852 43002
rect 7864 42950 7916 43002
rect 12047 42950 12099 43002
rect 12111 42950 12163 43002
rect 12175 42950 12227 43002
rect 12239 42950 12291 43002
rect 12303 42950 12355 43002
rect 16486 42950 16538 43002
rect 16550 42950 16602 43002
rect 16614 42950 16666 43002
rect 16678 42950 16730 43002
rect 16742 42950 16794 43002
rect 5388 42406 5440 42458
rect 5452 42406 5504 42458
rect 5516 42406 5568 42458
rect 5580 42406 5632 42458
rect 5644 42406 5696 42458
rect 9827 42406 9879 42458
rect 9891 42406 9943 42458
rect 9955 42406 10007 42458
rect 10019 42406 10071 42458
rect 10083 42406 10135 42458
rect 14266 42406 14318 42458
rect 14330 42406 14382 42458
rect 14394 42406 14446 42458
rect 14458 42406 14510 42458
rect 14522 42406 14574 42458
rect 18705 42406 18757 42458
rect 18769 42406 18821 42458
rect 18833 42406 18885 42458
rect 18897 42406 18949 42458
rect 18961 42406 19013 42458
rect 3169 41862 3221 41914
rect 3233 41862 3285 41914
rect 3297 41862 3349 41914
rect 3361 41862 3413 41914
rect 3425 41862 3477 41914
rect 7608 41862 7660 41914
rect 7672 41862 7724 41914
rect 7736 41862 7788 41914
rect 7800 41862 7852 41914
rect 7864 41862 7916 41914
rect 12047 41862 12099 41914
rect 12111 41862 12163 41914
rect 12175 41862 12227 41914
rect 12239 41862 12291 41914
rect 12303 41862 12355 41914
rect 16486 41862 16538 41914
rect 16550 41862 16602 41914
rect 16614 41862 16666 41914
rect 16678 41862 16730 41914
rect 16742 41862 16794 41914
rect 5388 41318 5440 41370
rect 5452 41318 5504 41370
rect 5516 41318 5568 41370
rect 5580 41318 5632 41370
rect 5644 41318 5696 41370
rect 9827 41318 9879 41370
rect 9891 41318 9943 41370
rect 9955 41318 10007 41370
rect 10019 41318 10071 41370
rect 10083 41318 10135 41370
rect 14266 41318 14318 41370
rect 14330 41318 14382 41370
rect 14394 41318 14446 41370
rect 14458 41318 14510 41370
rect 14522 41318 14574 41370
rect 18705 41318 18757 41370
rect 18769 41318 18821 41370
rect 18833 41318 18885 41370
rect 18897 41318 18949 41370
rect 18961 41318 19013 41370
rect 18328 41123 18380 41132
rect 18328 41089 18337 41123
rect 18337 41089 18371 41123
rect 18371 41089 18380 41123
rect 18328 41080 18380 41089
rect 18052 41012 18104 41064
rect 3169 40774 3221 40826
rect 3233 40774 3285 40826
rect 3297 40774 3349 40826
rect 3361 40774 3413 40826
rect 3425 40774 3477 40826
rect 7608 40774 7660 40826
rect 7672 40774 7724 40826
rect 7736 40774 7788 40826
rect 7800 40774 7852 40826
rect 7864 40774 7916 40826
rect 12047 40774 12099 40826
rect 12111 40774 12163 40826
rect 12175 40774 12227 40826
rect 12239 40774 12291 40826
rect 12303 40774 12355 40826
rect 16486 40774 16538 40826
rect 16550 40774 16602 40826
rect 16614 40774 16666 40826
rect 16678 40774 16730 40826
rect 16742 40774 16794 40826
rect 18328 40332 18380 40384
rect 5388 40230 5440 40282
rect 5452 40230 5504 40282
rect 5516 40230 5568 40282
rect 5580 40230 5632 40282
rect 5644 40230 5696 40282
rect 9827 40230 9879 40282
rect 9891 40230 9943 40282
rect 9955 40230 10007 40282
rect 10019 40230 10071 40282
rect 10083 40230 10135 40282
rect 14266 40230 14318 40282
rect 14330 40230 14382 40282
rect 14394 40230 14446 40282
rect 14458 40230 14510 40282
rect 14522 40230 14574 40282
rect 18705 40230 18757 40282
rect 18769 40230 18821 40282
rect 18833 40230 18885 40282
rect 18897 40230 18949 40282
rect 18961 40230 19013 40282
rect 3169 39686 3221 39738
rect 3233 39686 3285 39738
rect 3297 39686 3349 39738
rect 3361 39686 3413 39738
rect 3425 39686 3477 39738
rect 7608 39686 7660 39738
rect 7672 39686 7724 39738
rect 7736 39686 7788 39738
rect 7800 39686 7852 39738
rect 7864 39686 7916 39738
rect 12047 39686 12099 39738
rect 12111 39686 12163 39738
rect 12175 39686 12227 39738
rect 12239 39686 12291 39738
rect 12303 39686 12355 39738
rect 16486 39686 16538 39738
rect 16550 39686 16602 39738
rect 16614 39686 16666 39738
rect 16678 39686 16730 39738
rect 16742 39686 16794 39738
rect 5388 39142 5440 39194
rect 5452 39142 5504 39194
rect 5516 39142 5568 39194
rect 5580 39142 5632 39194
rect 5644 39142 5696 39194
rect 9827 39142 9879 39194
rect 9891 39142 9943 39194
rect 9955 39142 10007 39194
rect 10019 39142 10071 39194
rect 10083 39142 10135 39194
rect 14266 39142 14318 39194
rect 14330 39142 14382 39194
rect 14394 39142 14446 39194
rect 14458 39142 14510 39194
rect 14522 39142 14574 39194
rect 18705 39142 18757 39194
rect 18769 39142 18821 39194
rect 18833 39142 18885 39194
rect 18897 39142 18949 39194
rect 18961 39142 19013 39194
rect 3169 38598 3221 38650
rect 3233 38598 3285 38650
rect 3297 38598 3349 38650
rect 3361 38598 3413 38650
rect 3425 38598 3477 38650
rect 7608 38598 7660 38650
rect 7672 38598 7724 38650
rect 7736 38598 7788 38650
rect 7800 38598 7852 38650
rect 7864 38598 7916 38650
rect 12047 38598 12099 38650
rect 12111 38598 12163 38650
rect 12175 38598 12227 38650
rect 12239 38598 12291 38650
rect 12303 38598 12355 38650
rect 16486 38598 16538 38650
rect 16550 38598 16602 38650
rect 16614 38598 16666 38650
rect 16678 38598 16730 38650
rect 16742 38598 16794 38650
rect 5388 38054 5440 38106
rect 5452 38054 5504 38106
rect 5516 38054 5568 38106
rect 5580 38054 5632 38106
rect 5644 38054 5696 38106
rect 9827 38054 9879 38106
rect 9891 38054 9943 38106
rect 9955 38054 10007 38106
rect 10019 38054 10071 38106
rect 10083 38054 10135 38106
rect 14266 38054 14318 38106
rect 14330 38054 14382 38106
rect 14394 38054 14446 38106
rect 14458 38054 14510 38106
rect 14522 38054 14574 38106
rect 18705 38054 18757 38106
rect 18769 38054 18821 38106
rect 18833 38054 18885 38106
rect 18897 38054 18949 38106
rect 18961 38054 19013 38106
rect 3169 37510 3221 37562
rect 3233 37510 3285 37562
rect 3297 37510 3349 37562
rect 3361 37510 3413 37562
rect 3425 37510 3477 37562
rect 7608 37510 7660 37562
rect 7672 37510 7724 37562
rect 7736 37510 7788 37562
rect 7800 37510 7852 37562
rect 7864 37510 7916 37562
rect 12047 37510 12099 37562
rect 12111 37510 12163 37562
rect 12175 37510 12227 37562
rect 12239 37510 12291 37562
rect 12303 37510 12355 37562
rect 16486 37510 16538 37562
rect 16550 37510 16602 37562
rect 16614 37510 16666 37562
rect 16678 37510 16730 37562
rect 16742 37510 16794 37562
rect 5388 36966 5440 37018
rect 5452 36966 5504 37018
rect 5516 36966 5568 37018
rect 5580 36966 5632 37018
rect 5644 36966 5696 37018
rect 9827 36966 9879 37018
rect 9891 36966 9943 37018
rect 9955 36966 10007 37018
rect 10019 36966 10071 37018
rect 10083 36966 10135 37018
rect 14266 36966 14318 37018
rect 14330 36966 14382 37018
rect 14394 36966 14446 37018
rect 14458 36966 14510 37018
rect 14522 36966 14574 37018
rect 18705 36966 18757 37018
rect 18769 36966 18821 37018
rect 18833 36966 18885 37018
rect 18897 36966 18949 37018
rect 18961 36966 19013 37018
rect 3169 36422 3221 36474
rect 3233 36422 3285 36474
rect 3297 36422 3349 36474
rect 3361 36422 3413 36474
rect 3425 36422 3477 36474
rect 7608 36422 7660 36474
rect 7672 36422 7724 36474
rect 7736 36422 7788 36474
rect 7800 36422 7852 36474
rect 7864 36422 7916 36474
rect 12047 36422 12099 36474
rect 12111 36422 12163 36474
rect 12175 36422 12227 36474
rect 12239 36422 12291 36474
rect 12303 36422 12355 36474
rect 16486 36422 16538 36474
rect 16550 36422 16602 36474
rect 16614 36422 16666 36474
rect 16678 36422 16730 36474
rect 16742 36422 16794 36474
rect 5388 35878 5440 35930
rect 5452 35878 5504 35930
rect 5516 35878 5568 35930
rect 5580 35878 5632 35930
rect 5644 35878 5696 35930
rect 9827 35878 9879 35930
rect 9891 35878 9943 35930
rect 9955 35878 10007 35930
rect 10019 35878 10071 35930
rect 10083 35878 10135 35930
rect 14266 35878 14318 35930
rect 14330 35878 14382 35930
rect 14394 35878 14446 35930
rect 14458 35878 14510 35930
rect 14522 35878 14574 35930
rect 18705 35878 18757 35930
rect 18769 35878 18821 35930
rect 18833 35878 18885 35930
rect 18897 35878 18949 35930
rect 18961 35878 19013 35930
rect 3169 35334 3221 35386
rect 3233 35334 3285 35386
rect 3297 35334 3349 35386
rect 3361 35334 3413 35386
rect 3425 35334 3477 35386
rect 7608 35334 7660 35386
rect 7672 35334 7724 35386
rect 7736 35334 7788 35386
rect 7800 35334 7852 35386
rect 7864 35334 7916 35386
rect 12047 35334 12099 35386
rect 12111 35334 12163 35386
rect 12175 35334 12227 35386
rect 12239 35334 12291 35386
rect 12303 35334 12355 35386
rect 16486 35334 16538 35386
rect 16550 35334 16602 35386
rect 16614 35334 16666 35386
rect 16678 35334 16730 35386
rect 16742 35334 16794 35386
rect 5388 34790 5440 34842
rect 5452 34790 5504 34842
rect 5516 34790 5568 34842
rect 5580 34790 5632 34842
rect 5644 34790 5696 34842
rect 9827 34790 9879 34842
rect 9891 34790 9943 34842
rect 9955 34790 10007 34842
rect 10019 34790 10071 34842
rect 10083 34790 10135 34842
rect 14266 34790 14318 34842
rect 14330 34790 14382 34842
rect 14394 34790 14446 34842
rect 14458 34790 14510 34842
rect 14522 34790 14574 34842
rect 18705 34790 18757 34842
rect 18769 34790 18821 34842
rect 18833 34790 18885 34842
rect 18897 34790 18949 34842
rect 18961 34790 19013 34842
rect 18512 34391 18564 34400
rect 18512 34357 18521 34391
rect 18521 34357 18555 34391
rect 18555 34357 18564 34391
rect 18512 34348 18564 34357
rect 3169 34246 3221 34298
rect 3233 34246 3285 34298
rect 3297 34246 3349 34298
rect 3361 34246 3413 34298
rect 3425 34246 3477 34298
rect 7608 34246 7660 34298
rect 7672 34246 7724 34298
rect 7736 34246 7788 34298
rect 7800 34246 7852 34298
rect 7864 34246 7916 34298
rect 12047 34246 12099 34298
rect 12111 34246 12163 34298
rect 12175 34246 12227 34298
rect 12239 34246 12291 34298
rect 12303 34246 12355 34298
rect 16486 34246 16538 34298
rect 16550 34246 16602 34298
rect 16614 34246 16666 34298
rect 16678 34246 16730 34298
rect 16742 34246 16794 34298
rect 5388 33702 5440 33754
rect 5452 33702 5504 33754
rect 5516 33702 5568 33754
rect 5580 33702 5632 33754
rect 5644 33702 5696 33754
rect 9827 33702 9879 33754
rect 9891 33702 9943 33754
rect 9955 33702 10007 33754
rect 10019 33702 10071 33754
rect 10083 33702 10135 33754
rect 14266 33702 14318 33754
rect 14330 33702 14382 33754
rect 14394 33702 14446 33754
rect 14458 33702 14510 33754
rect 14522 33702 14574 33754
rect 18705 33702 18757 33754
rect 18769 33702 18821 33754
rect 18833 33702 18885 33754
rect 18897 33702 18949 33754
rect 18961 33702 19013 33754
rect 3169 33158 3221 33210
rect 3233 33158 3285 33210
rect 3297 33158 3349 33210
rect 3361 33158 3413 33210
rect 3425 33158 3477 33210
rect 7608 33158 7660 33210
rect 7672 33158 7724 33210
rect 7736 33158 7788 33210
rect 7800 33158 7852 33210
rect 7864 33158 7916 33210
rect 12047 33158 12099 33210
rect 12111 33158 12163 33210
rect 12175 33158 12227 33210
rect 12239 33158 12291 33210
rect 12303 33158 12355 33210
rect 16486 33158 16538 33210
rect 16550 33158 16602 33210
rect 16614 33158 16666 33210
rect 16678 33158 16730 33210
rect 16742 33158 16794 33210
rect 5388 32614 5440 32666
rect 5452 32614 5504 32666
rect 5516 32614 5568 32666
rect 5580 32614 5632 32666
rect 5644 32614 5696 32666
rect 9827 32614 9879 32666
rect 9891 32614 9943 32666
rect 9955 32614 10007 32666
rect 10019 32614 10071 32666
rect 10083 32614 10135 32666
rect 14266 32614 14318 32666
rect 14330 32614 14382 32666
rect 14394 32614 14446 32666
rect 14458 32614 14510 32666
rect 14522 32614 14574 32666
rect 18705 32614 18757 32666
rect 18769 32614 18821 32666
rect 18833 32614 18885 32666
rect 18897 32614 18949 32666
rect 18961 32614 19013 32666
rect 3169 32070 3221 32122
rect 3233 32070 3285 32122
rect 3297 32070 3349 32122
rect 3361 32070 3413 32122
rect 3425 32070 3477 32122
rect 7608 32070 7660 32122
rect 7672 32070 7724 32122
rect 7736 32070 7788 32122
rect 7800 32070 7852 32122
rect 7864 32070 7916 32122
rect 12047 32070 12099 32122
rect 12111 32070 12163 32122
rect 12175 32070 12227 32122
rect 12239 32070 12291 32122
rect 12303 32070 12355 32122
rect 16486 32070 16538 32122
rect 16550 32070 16602 32122
rect 16614 32070 16666 32122
rect 16678 32070 16730 32122
rect 16742 32070 16794 32122
rect 5388 31526 5440 31578
rect 5452 31526 5504 31578
rect 5516 31526 5568 31578
rect 5580 31526 5632 31578
rect 5644 31526 5696 31578
rect 9827 31526 9879 31578
rect 9891 31526 9943 31578
rect 9955 31526 10007 31578
rect 10019 31526 10071 31578
rect 10083 31526 10135 31578
rect 14266 31526 14318 31578
rect 14330 31526 14382 31578
rect 14394 31526 14446 31578
rect 14458 31526 14510 31578
rect 14522 31526 14574 31578
rect 18705 31526 18757 31578
rect 18769 31526 18821 31578
rect 18833 31526 18885 31578
rect 18897 31526 18949 31578
rect 18961 31526 19013 31578
rect 3169 30982 3221 31034
rect 3233 30982 3285 31034
rect 3297 30982 3349 31034
rect 3361 30982 3413 31034
rect 3425 30982 3477 31034
rect 7608 30982 7660 31034
rect 7672 30982 7724 31034
rect 7736 30982 7788 31034
rect 7800 30982 7852 31034
rect 7864 30982 7916 31034
rect 12047 30982 12099 31034
rect 12111 30982 12163 31034
rect 12175 30982 12227 31034
rect 12239 30982 12291 31034
rect 12303 30982 12355 31034
rect 16486 30982 16538 31034
rect 16550 30982 16602 31034
rect 16614 30982 16666 31034
rect 16678 30982 16730 31034
rect 16742 30982 16794 31034
rect 5388 30438 5440 30490
rect 5452 30438 5504 30490
rect 5516 30438 5568 30490
rect 5580 30438 5632 30490
rect 5644 30438 5696 30490
rect 9827 30438 9879 30490
rect 9891 30438 9943 30490
rect 9955 30438 10007 30490
rect 10019 30438 10071 30490
rect 10083 30438 10135 30490
rect 14266 30438 14318 30490
rect 14330 30438 14382 30490
rect 14394 30438 14446 30490
rect 14458 30438 14510 30490
rect 14522 30438 14574 30490
rect 18705 30438 18757 30490
rect 18769 30438 18821 30490
rect 18833 30438 18885 30490
rect 18897 30438 18949 30490
rect 18961 30438 19013 30490
rect 3169 29894 3221 29946
rect 3233 29894 3285 29946
rect 3297 29894 3349 29946
rect 3361 29894 3413 29946
rect 3425 29894 3477 29946
rect 7608 29894 7660 29946
rect 7672 29894 7724 29946
rect 7736 29894 7788 29946
rect 7800 29894 7852 29946
rect 7864 29894 7916 29946
rect 12047 29894 12099 29946
rect 12111 29894 12163 29946
rect 12175 29894 12227 29946
rect 12239 29894 12291 29946
rect 12303 29894 12355 29946
rect 16486 29894 16538 29946
rect 16550 29894 16602 29946
rect 16614 29894 16666 29946
rect 16678 29894 16730 29946
rect 16742 29894 16794 29946
rect 5388 29350 5440 29402
rect 5452 29350 5504 29402
rect 5516 29350 5568 29402
rect 5580 29350 5632 29402
rect 5644 29350 5696 29402
rect 9827 29350 9879 29402
rect 9891 29350 9943 29402
rect 9955 29350 10007 29402
rect 10019 29350 10071 29402
rect 10083 29350 10135 29402
rect 14266 29350 14318 29402
rect 14330 29350 14382 29402
rect 14394 29350 14446 29402
rect 14458 29350 14510 29402
rect 14522 29350 14574 29402
rect 18705 29350 18757 29402
rect 18769 29350 18821 29402
rect 18833 29350 18885 29402
rect 18897 29350 18949 29402
rect 18961 29350 19013 29402
rect 3169 28806 3221 28858
rect 3233 28806 3285 28858
rect 3297 28806 3349 28858
rect 3361 28806 3413 28858
rect 3425 28806 3477 28858
rect 7608 28806 7660 28858
rect 7672 28806 7724 28858
rect 7736 28806 7788 28858
rect 7800 28806 7852 28858
rect 7864 28806 7916 28858
rect 12047 28806 12099 28858
rect 12111 28806 12163 28858
rect 12175 28806 12227 28858
rect 12239 28806 12291 28858
rect 12303 28806 12355 28858
rect 16486 28806 16538 28858
rect 16550 28806 16602 28858
rect 16614 28806 16666 28858
rect 16678 28806 16730 28858
rect 16742 28806 16794 28858
rect 18604 28432 18656 28484
rect 17040 28407 17092 28416
rect 17040 28373 17049 28407
rect 17049 28373 17083 28407
rect 17083 28373 17092 28407
rect 17040 28364 17092 28373
rect 5388 28262 5440 28314
rect 5452 28262 5504 28314
rect 5516 28262 5568 28314
rect 5580 28262 5632 28314
rect 5644 28262 5696 28314
rect 9827 28262 9879 28314
rect 9891 28262 9943 28314
rect 9955 28262 10007 28314
rect 10019 28262 10071 28314
rect 10083 28262 10135 28314
rect 14266 28262 14318 28314
rect 14330 28262 14382 28314
rect 14394 28262 14446 28314
rect 14458 28262 14510 28314
rect 14522 28262 14574 28314
rect 18705 28262 18757 28314
rect 18769 28262 18821 28314
rect 18833 28262 18885 28314
rect 18897 28262 18949 28314
rect 18961 28262 19013 28314
rect 3169 27718 3221 27770
rect 3233 27718 3285 27770
rect 3297 27718 3349 27770
rect 3361 27718 3413 27770
rect 3425 27718 3477 27770
rect 7608 27718 7660 27770
rect 7672 27718 7724 27770
rect 7736 27718 7788 27770
rect 7800 27718 7852 27770
rect 7864 27718 7916 27770
rect 12047 27718 12099 27770
rect 12111 27718 12163 27770
rect 12175 27718 12227 27770
rect 12239 27718 12291 27770
rect 12303 27718 12355 27770
rect 16486 27718 16538 27770
rect 16550 27718 16602 27770
rect 16614 27718 16666 27770
rect 16678 27718 16730 27770
rect 16742 27718 16794 27770
rect 5388 27174 5440 27226
rect 5452 27174 5504 27226
rect 5516 27174 5568 27226
rect 5580 27174 5632 27226
rect 5644 27174 5696 27226
rect 9827 27174 9879 27226
rect 9891 27174 9943 27226
rect 9955 27174 10007 27226
rect 10019 27174 10071 27226
rect 10083 27174 10135 27226
rect 14266 27174 14318 27226
rect 14330 27174 14382 27226
rect 14394 27174 14446 27226
rect 14458 27174 14510 27226
rect 14522 27174 14574 27226
rect 18705 27174 18757 27226
rect 18769 27174 18821 27226
rect 18833 27174 18885 27226
rect 18897 27174 18949 27226
rect 18961 27174 19013 27226
rect 3169 26630 3221 26682
rect 3233 26630 3285 26682
rect 3297 26630 3349 26682
rect 3361 26630 3413 26682
rect 3425 26630 3477 26682
rect 7608 26630 7660 26682
rect 7672 26630 7724 26682
rect 7736 26630 7788 26682
rect 7800 26630 7852 26682
rect 7864 26630 7916 26682
rect 12047 26630 12099 26682
rect 12111 26630 12163 26682
rect 12175 26630 12227 26682
rect 12239 26630 12291 26682
rect 12303 26630 12355 26682
rect 16486 26630 16538 26682
rect 16550 26630 16602 26682
rect 16614 26630 16666 26682
rect 16678 26630 16730 26682
rect 16742 26630 16794 26682
rect 5388 26086 5440 26138
rect 5452 26086 5504 26138
rect 5516 26086 5568 26138
rect 5580 26086 5632 26138
rect 5644 26086 5696 26138
rect 9827 26086 9879 26138
rect 9891 26086 9943 26138
rect 9955 26086 10007 26138
rect 10019 26086 10071 26138
rect 10083 26086 10135 26138
rect 14266 26086 14318 26138
rect 14330 26086 14382 26138
rect 14394 26086 14446 26138
rect 14458 26086 14510 26138
rect 14522 26086 14574 26138
rect 18705 26086 18757 26138
rect 18769 26086 18821 26138
rect 18833 26086 18885 26138
rect 18897 26086 18949 26138
rect 18961 26086 19013 26138
rect 3169 25542 3221 25594
rect 3233 25542 3285 25594
rect 3297 25542 3349 25594
rect 3361 25542 3413 25594
rect 3425 25542 3477 25594
rect 7608 25542 7660 25594
rect 7672 25542 7724 25594
rect 7736 25542 7788 25594
rect 7800 25542 7852 25594
rect 7864 25542 7916 25594
rect 12047 25542 12099 25594
rect 12111 25542 12163 25594
rect 12175 25542 12227 25594
rect 12239 25542 12291 25594
rect 12303 25542 12355 25594
rect 16486 25542 16538 25594
rect 16550 25542 16602 25594
rect 16614 25542 16666 25594
rect 16678 25542 16730 25594
rect 16742 25542 16794 25594
rect 5388 24998 5440 25050
rect 5452 24998 5504 25050
rect 5516 24998 5568 25050
rect 5580 24998 5632 25050
rect 5644 24998 5696 25050
rect 9827 24998 9879 25050
rect 9891 24998 9943 25050
rect 9955 24998 10007 25050
rect 10019 24998 10071 25050
rect 10083 24998 10135 25050
rect 14266 24998 14318 25050
rect 14330 24998 14382 25050
rect 14394 24998 14446 25050
rect 14458 24998 14510 25050
rect 14522 24998 14574 25050
rect 18705 24998 18757 25050
rect 18769 24998 18821 25050
rect 18833 24998 18885 25050
rect 18897 24998 18949 25050
rect 18961 24998 19013 25050
rect 3169 24454 3221 24506
rect 3233 24454 3285 24506
rect 3297 24454 3349 24506
rect 3361 24454 3413 24506
rect 3425 24454 3477 24506
rect 7608 24454 7660 24506
rect 7672 24454 7724 24506
rect 7736 24454 7788 24506
rect 7800 24454 7852 24506
rect 7864 24454 7916 24506
rect 12047 24454 12099 24506
rect 12111 24454 12163 24506
rect 12175 24454 12227 24506
rect 12239 24454 12291 24506
rect 12303 24454 12355 24506
rect 16486 24454 16538 24506
rect 16550 24454 16602 24506
rect 16614 24454 16666 24506
rect 16678 24454 16730 24506
rect 16742 24454 16794 24506
rect 5388 23910 5440 23962
rect 5452 23910 5504 23962
rect 5516 23910 5568 23962
rect 5580 23910 5632 23962
rect 5644 23910 5696 23962
rect 9827 23910 9879 23962
rect 9891 23910 9943 23962
rect 9955 23910 10007 23962
rect 10019 23910 10071 23962
rect 10083 23910 10135 23962
rect 14266 23910 14318 23962
rect 14330 23910 14382 23962
rect 14394 23910 14446 23962
rect 14458 23910 14510 23962
rect 14522 23910 14574 23962
rect 18705 23910 18757 23962
rect 18769 23910 18821 23962
rect 18833 23910 18885 23962
rect 18897 23910 18949 23962
rect 18961 23910 19013 23962
rect 3169 23366 3221 23418
rect 3233 23366 3285 23418
rect 3297 23366 3349 23418
rect 3361 23366 3413 23418
rect 3425 23366 3477 23418
rect 7608 23366 7660 23418
rect 7672 23366 7724 23418
rect 7736 23366 7788 23418
rect 7800 23366 7852 23418
rect 7864 23366 7916 23418
rect 12047 23366 12099 23418
rect 12111 23366 12163 23418
rect 12175 23366 12227 23418
rect 12239 23366 12291 23418
rect 12303 23366 12355 23418
rect 16486 23366 16538 23418
rect 16550 23366 16602 23418
rect 16614 23366 16666 23418
rect 16678 23366 16730 23418
rect 16742 23366 16794 23418
rect 5388 22822 5440 22874
rect 5452 22822 5504 22874
rect 5516 22822 5568 22874
rect 5580 22822 5632 22874
rect 5644 22822 5696 22874
rect 9827 22822 9879 22874
rect 9891 22822 9943 22874
rect 9955 22822 10007 22874
rect 10019 22822 10071 22874
rect 10083 22822 10135 22874
rect 14266 22822 14318 22874
rect 14330 22822 14382 22874
rect 14394 22822 14446 22874
rect 14458 22822 14510 22874
rect 14522 22822 14574 22874
rect 18705 22822 18757 22874
rect 18769 22822 18821 22874
rect 18833 22822 18885 22874
rect 18897 22822 18949 22874
rect 18961 22822 19013 22874
rect 3169 22278 3221 22330
rect 3233 22278 3285 22330
rect 3297 22278 3349 22330
rect 3361 22278 3413 22330
rect 3425 22278 3477 22330
rect 7608 22278 7660 22330
rect 7672 22278 7724 22330
rect 7736 22278 7788 22330
rect 7800 22278 7852 22330
rect 7864 22278 7916 22330
rect 12047 22278 12099 22330
rect 12111 22278 12163 22330
rect 12175 22278 12227 22330
rect 12239 22278 12291 22330
rect 12303 22278 12355 22330
rect 16486 22278 16538 22330
rect 16550 22278 16602 22330
rect 16614 22278 16666 22330
rect 16678 22278 16730 22330
rect 16742 22278 16794 22330
rect 18512 22219 18564 22228
rect 18512 22185 18521 22219
rect 18521 22185 18555 22219
rect 18555 22185 18564 22219
rect 18512 22176 18564 22185
rect 5388 21734 5440 21786
rect 5452 21734 5504 21786
rect 5516 21734 5568 21786
rect 5580 21734 5632 21786
rect 5644 21734 5696 21786
rect 9827 21734 9879 21786
rect 9891 21734 9943 21786
rect 9955 21734 10007 21786
rect 10019 21734 10071 21786
rect 10083 21734 10135 21786
rect 14266 21734 14318 21786
rect 14330 21734 14382 21786
rect 14394 21734 14446 21786
rect 14458 21734 14510 21786
rect 14522 21734 14574 21786
rect 18705 21734 18757 21786
rect 18769 21734 18821 21786
rect 18833 21734 18885 21786
rect 18897 21734 18949 21786
rect 18961 21734 19013 21786
rect 3169 21190 3221 21242
rect 3233 21190 3285 21242
rect 3297 21190 3349 21242
rect 3361 21190 3413 21242
rect 3425 21190 3477 21242
rect 7608 21190 7660 21242
rect 7672 21190 7724 21242
rect 7736 21190 7788 21242
rect 7800 21190 7852 21242
rect 7864 21190 7916 21242
rect 12047 21190 12099 21242
rect 12111 21190 12163 21242
rect 12175 21190 12227 21242
rect 12239 21190 12291 21242
rect 12303 21190 12355 21242
rect 16486 21190 16538 21242
rect 16550 21190 16602 21242
rect 16614 21190 16666 21242
rect 16678 21190 16730 21242
rect 16742 21190 16794 21242
rect 5388 20646 5440 20698
rect 5452 20646 5504 20698
rect 5516 20646 5568 20698
rect 5580 20646 5632 20698
rect 5644 20646 5696 20698
rect 9827 20646 9879 20698
rect 9891 20646 9943 20698
rect 9955 20646 10007 20698
rect 10019 20646 10071 20698
rect 10083 20646 10135 20698
rect 14266 20646 14318 20698
rect 14330 20646 14382 20698
rect 14394 20646 14446 20698
rect 14458 20646 14510 20698
rect 14522 20646 14574 20698
rect 18705 20646 18757 20698
rect 18769 20646 18821 20698
rect 18833 20646 18885 20698
rect 18897 20646 18949 20698
rect 18961 20646 19013 20698
rect 3169 20102 3221 20154
rect 3233 20102 3285 20154
rect 3297 20102 3349 20154
rect 3361 20102 3413 20154
rect 3425 20102 3477 20154
rect 7608 20102 7660 20154
rect 7672 20102 7724 20154
rect 7736 20102 7788 20154
rect 7800 20102 7852 20154
rect 7864 20102 7916 20154
rect 12047 20102 12099 20154
rect 12111 20102 12163 20154
rect 12175 20102 12227 20154
rect 12239 20102 12291 20154
rect 12303 20102 12355 20154
rect 16486 20102 16538 20154
rect 16550 20102 16602 20154
rect 16614 20102 16666 20154
rect 16678 20102 16730 20154
rect 16742 20102 16794 20154
rect 5388 19558 5440 19610
rect 5452 19558 5504 19610
rect 5516 19558 5568 19610
rect 5580 19558 5632 19610
rect 5644 19558 5696 19610
rect 9827 19558 9879 19610
rect 9891 19558 9943 19610
rect 9955 19558 10007 19610
rect 10019 19558 10071 19610
rect 10083 19558 10135 19610
rect 14266 19558 14318 19610
rect 14330 19558 14382 19610
rect 14394 19558 14446 19610
rect 14458 19558 14510 19610
rect 14522 19558 14574 19610
rect 18705 19558 18757 19610
rect 18769 19558 18821 19610
rect 18833 19558 18885 19610
rect 18897 19558 18949 19610
rect 18961 19558 19013 19610
rect 3169 19014 3221 19066
rect 3233 19014 3285 19066
rect 3297 19014 3349 19066
rect 3361 19014 3413 19066
rect 3425 19014 3477 19066
rect 7608 19014 7660 19066
rect 7672 19014 7724 19066
rect 7736 19014 7788 19066
rect 7800 19014 7852 19066
rect 7864 19014 7916 19066
rect 12047 19014 12099 19066
rect 12111 19014 12163 19066
rect 12175 19014 12227 19066
rect 12239 19014 12291 19066
rect 12303 19014 12355 19066
rect 16486 19014 16538 19066
rect 16550 19014 16602 19066
rect 16614 19014 16666 19066
rect 16678 19014 16730 19066
rect 16742 19014 16794 19066
rect 5388 18470 5440 18522
rect 5452 18470 5504 18522
rect 5516 18470 5568 18522
rect 5580 18470 5632 18522
rect 5644 18470 5696 18522
rect 9827 18470 9879 18522
rect 9891 18470 9943 18522
rect 9955 18470 10007 18522
rect 10019 18470 10071 18522
rect 10083 18470 10135 18522
rect 14266 18470 14318 18522
rect 14330 18470 14382 18522
rect 14394 18470 14446 18522
rect 14458 18470 14510 18522
rect 14522 18470 14574 18522
rect 18705 18470 18757 18522
rect 18769 18470 18821 18522
rect 18833 18470 18885 18522
rect 18897 18470 18949 18522
rect 18961 18470 19013 18522
rect 3169 17926 3221 17978
rect 3233 17926 3285 17978
rect 3297 17926 3349 17978
rect 3361 17926 3413 17978
rect 3425 17926 3477 17978
rect 7608 17926 7660 17978
rect 7672 17926 7724 17978
rect 7736 17926 7788 17978
rect 7800 17926 7852 17978
rect 7864 17926 7916 17978
rect 12047 17926 12099 17978
rect 12111 17926 12163 17978
rect 12175 17926 12227 17978
rect 12239 17926 12291 17978
rect 12303 17926 12355 17978
rect 16486 17926 16538 17978
rect 16550 17926 16602 17978
rect 16614 17926 16666 17978
rect 16678 17926 16730 17978
rect 16742 17926 16794 17978
rect 5388 17382 5440 17434
rect 5452 17382 5504 17434
rect 5516 17382 5568 17434
rect 5580 17382 5632 17434
rect 5644 17382 5696 17434
rect 9827 17382 9879 17434
rect 9891 17382 9943 17434
rect 9955 17382 10007 17434
rect 10019 17382 10071 17434
rect 10083 17382 10135 17434
rect 14266 17382 14318 17434
rect 14330 17382 14382 17434
rect 14394 17382 14446 17434
rect 14458 17382 14510 17434
rect 14522 17382 14574 17434
rect 18705 17382 18757 17434
rect 18769 17382 18821 17434
rect 18833 17382 18885 17434
rect 18897 17382 18949 17434
rect 18961 17382 19013 17434
rect 3169 16838 3221 16890
rect 3233 16838 3285 16890
rect 3297 16838 3349 16890
rect 3361 16838 3413 16890
rect 3425 16838 3477 16890
rect 7608 16838 7660 16890
rect 7672 16838 7724 16890
rect 7736 16838 7788 16890
rect 7800 16838 7852 16890
rect 7864 16838 7916 16890
rect 12047 16838 12099 16890
rect 12111 16838 12163 16890
rect 12175 16838 12227 16890
rect 12239 16838 12291 16890
rect 12303 16838 12355 16890
rect 16486 16838 16538 16890
rect 16550 16838 16602 16890
rect 16614 16838 16666 16890
rect 16678 16838 16730 16890
rect 16742 16838 16794 16890
rect 5388 16294 5440 16346
rect 5452 16294 5504 16346
rect 5516 16294 5568 16346
rect 5580 16294 5632 16346
rect 5644 16294 5696 16346
rect 9827 16294 9879 16346
rect 9891 16294 9943 16346
rect 9955 16294 10007 16346
rect 10019 16294 10071 16346
rect 10083 16294 10135 16346
rect 14266 16294 14318 16346
rect 14330 16294 14382 16346
rect 14394 16294 14446 16346
rect 14458 16294 14510 16346
rect 14522 16294 14574 16346
rect 18705 16294 18757 16346
rect 18769 16294 18821 16346
rect 18833 16294 18885 16346
rect 18897 16294 18949 16346
rect 18961 16294 19013 16346
rect 17132 16099 17184 16108
rect 17132 16065 17141 16099
rect 17141 16065 17175 16099
rect 17175 16065 17184 16099
rect 17132 16056 17184 16065
rect 18328 16031 18380 16040
rect 18328 15997 18337 16031
rect 18337 15997 18371 16031
rect 18371 15997 18380 16031
rect 18328 15988 18380 15997
rect 3169 15750 3221 15802
rect 3233 15750 3285 15802
rect 3297 15750 3349 15802
rect 3361 15750 3413 15802
rect 3425 15750 3477 15802
rect 7608 15750 7660 15802
rect 7672 15750 7724 15802
rect 7736 15750 7788 15802
rect 7800 15750 7852 15802
rect 7864 15750 7916 15802
rect 12047 15750 12099 15802
rect 12111 15750 12163 15802
rect 12175 15750 12227 15802
rect 12239 15750 12291 15802
rect 12303 15750 12355 15802
rect 16486 15750 16538 15802
rect 16550 15750 16602 15802
rect 16614 15750 16666 15802
rect 16678 15750 16730 15802
rect 16742 15750 16794 15802
rect 5388 15206 5440 15258
rect 5452 15206 5504 15258
rect 5516 15206 5568 15258
rect 5580 15206 5632 15258
rect 5644 15206 5696 15258
rect 9827 15206 9879 15258
rect 9891 15206 9943 15258
rect 9955 15206 10007 15258
rect 10019 15206 10071 15258
rect 10083 15206 10135 15258
rect 14266 15206 14318 15258
rect 14330 15206 14382 15258
rect 14394 15206 14446 15258
rect 14458 15206 14510 15258
rect 14522 15206 14574 15258
rect 18705 15206 18757 15258
rect 18769 15206 18821 15258
rect 18833 15206 18885 15258
rect 18897 15206 18949 15258
rect 18961 15206 19013 15258
rect 3169 14662 3221 14714
rect 3233 14662 3285 14714
rect 3297 14662 3349 14714
rect 3361 14662 3413 14714
rect 3425 14662 3477 14714
rect 7608 14662 7660 14714
rect 7672 14662 7724 14714
rect 7736 14662 7788 14714
rect 7800 14662 7852 14714
rect 7864 14662 7916 14714
rect 12047 14662 12099 14714
rect 12111 14662 12163 14714
rect 12175 14662 12227 14714
rect 12239 14662 12291 14714
rect 12303 14662 12355 14714
rect 16486 14662 16538 14714
rect 16550 14662 16602 14714
rect 16614 14662 16666 14714
rect 16678 14662 16730 14714
rect 16742 14662 16794 14714
rect 5388 14118 5440 14170
rect 5452 14118 5504 14170
rect 5516 14118 5568 14170
rect 5580 14118 5632 14170
rect 5644 14118 5696 14170
rect 9827 14118 9879 14170
rect 9891 14118 9943 14170
rect 9955 14118 10007 14170
rect 10019 14118 10071 14170
rect 10083 14118 10135 14170
rect 14266 14118 14318 14170
rect 14330 14118 14382 14170
rect 14394 14118 14446 14170
rect 14458 14118 14510 14170
rect 14522 14118 14574 14170
rect 18705 14118 18757 14170
rect 18769 14118 18821 14170
rect 18833 14118 18885 14170
rect 18897 14118 18949 14170
rect 18961 14118 19013 14170
rect 3169 13574 3221 13626
rect 3233 13574 3285 13626
rect 3297 13574 3349 13626
rect 3361 13574 3413 13626
rect 3425 13574 3477 13626
rect 7608 13574 7660 13626
rect 7672 13574 7724 13626
rect 7736 13574 7788 13626
rect 7800 13574 7852 13626
rect 7864 13574 7916 13626
rect 12047 13574 12099 13626
rect 12111 13574 12163 13626
rect 12175 13574 12227 13626
rect 12239 13574 12291 13626
rect 12303 13574 12355 13626
rect 16486 13574 16538 13626
rect 16550 13574 16602 13626
rect 16614 13574 16666 13626
rect 16678 13574 16730 13626
rect 16742 13574 16794 13626
rect 5388 13030 5440 13082
rect 5452 13030 5504 13082
rect 5516 13030 5568 13082
rect 5580 13030 5632 13082
rect 5644 13030 5696 13082
rect 9827 13030 9879 13082
rect 9891 13030 9943 13082
rect 9955 13030 10007 13082
rect 10019 13030 10071 13082
rect 10083 13030 10135 13082
rect 14266 13030 14318 13082
rect 14330 13030 14382 13082
rect 14394 13030 14446 13082
rect 14458 13030 14510 13082
rect 14522 13030 14574 13082
rect 18705 13030 18757 13082
rect 18769 13030 18821 13082
rect 18833 13030 18885 13082
rect 18897 13030 18949 13082
rect 18961 13030 19013 13082
rect 3169 12486 3221 12538
rect 3233 12486 3285 12538
rect 3297 12486 3349 12538
rect 3361 12486 3413 12538
rect 3425 12486 3477 12538
rect 7608 12486 7660 12538
rect 7672 12486 7724 12538
rect 7736 12486 7788 12538
rect 7800 12486 7852 12538
rect 7864 12486 7916 12538
rect 12047 12486 12099 12538
rect 12111 12486 12163 12538
rect 12175 12486 12227 12538
rect 12239 12486 12291 12538
rect 12303 12486 12355 12538
rect 16486 12486 16538 12538
rect 16550 12486 16602 12538
rect 16614 12486 16666 12538
rect 16678 12486 16730 12538
rect 16742 12486 16794 12538
rect 5388 11942 5440 11994
rect 5452 11942 5504 11994
rect 5516 11942 5568 11994
rect 5580 11942 5632 11994
rect 5644 11942 5696 11994
rect 9827 11942 9879 11994
rect 9891 11942 9943 11994
rect 9955 11942 10007 11994
rect 10019 11942 10071 11994
rect 10083 11942 10135 11994
rect 14266 11942 14318 11994
rect 14330 11942 14382 11994
rect 14394 11942 14446 11994
rect 14458 11942 14510 11994
rect 14522 11942 14574 11994
rect 18705 11942 18757 11994
rect 18769 11942 18821 11994
rect 18833 11942 18885 11994
rect 18897 11942 18949 11994
rect 18961 11942 19013 11994
rect 3169 11398 3221 11450
rect 3233 11398 3285 11450
rect 3297 11398 3349 11450
rect 3361 11398 3413 11450
rect 3425 11398 3477 11450
rect 7608 11398 7660 11450
rect 7672 11398 7724 11450
rect 7736 11398 7788 11450
rect 7800 11398 7852 11450
rect 7864 11398 7916 11450
rect 12047 11398 12099 11450
rect 12111 11398 12163 11450
rect 12175 11398 12227 11450
rect 12239 11398 12291 11450
rect 12303 11398 12355 11450
rect 16486 11398 16538 11450
rect 16550 11398 16602 11450
rect 16614 11398 16666 11450
rect 16678 11398 16730 11450
rect 16742 11398 16794 11450
rect 5388 10854 5440 10906
rect 5452 10854 5504 10906
rect 5516 10854 5568 10906
rect 5580 10854 5632 10906
rect 5644 10854 5696 10906
rect 9827 10854 9879 10906
rect 9891 10854 9943 10906
rect 9955 10854 10007 10906
rect 10019 10854 10071 10906
rect 10083 10854 10135 10906
rect 14266 10854 14318 10906
rect 14330 10854 14382 10906
rect 14394 10854 14446 10906
rect 14458 10854 14510 10906
rect 14522 10854 14574 10906
rect 18705 10854 18757 10906
rect 18769 10854 18821 10906
rect 18833 10854 18885 10906
rect 18897 10854 18949 10906
rect 18961 10854 19013 10906
rect 3169 10310 3221 10362
rect 3233 10310 3285 10362
rect 3297 10310 3349 10362
rect 3361 10310 3413 10362
rect 3425 10310 3477 10362
rect 7608 10310 7660 10362
rect 7672 10310 7724 10362
rect 7736 10310 7788 10362
rect 7800 10310 7852 10362
rect 7864 10310 7916 10362
rect 12047 10310 12099 10362
rect 12111 10310 12163 10362
rect 12175 10310 12227 10362
rect 12239 10310 12291 10362
rect 12303 10310 12355 10362
rect 16486 10310 16538 10362
rect 16550 10310 16602 10362
rect 16614 10310 16666 10362
rect 16678 10310 16730 10362
rect 16742 10310 16794 10362
rect 5388 9766 5440 9818
rect 5452 9766 5504 9818
rect 5516 9766 5568 9818
rect 5580 9766 5632 9818
rect 5644 9766 5696 9818
rect 9827 9766 9879 9818
rect 9891 9766 9943 9818
rect 9955 9766 10007 9818
rect 10019 9766 10071 9818
rect 10083 9766 10135 9818
rect 14266 9766 14318 9818
rect 14330 9766 14382 9818
rect 14394 9766 14446 9818
rect 14458 9766 14510 9818
rect 14522 9766 14574 9818
rect 18705 9766 18757 9818
rect 18769 9766 18821 9818
rect 18833 9766 18885 9818
rect 18897 9766 18949 9818
rect 18961 9766 19013 9818
rect 18512 9367 18564 9376
rect 18512 9333 18521 9367
rect 18521 9333 18555 9367
rect 18555 9333 18564 9367
rect 18512 9324 18564 9333
rect 3169 9222 3221 9274
rect 3233 9222 3285 9274
rect 3297 9222 3349 9274
rect 3361 9222 3413 9274
rect 3425 9222 3477 9274
rect 7608 9222 7660 9274
rect 7672 9222 7724 9274
rect 7736 9222 7788 9274
rect 7800 9222 7852 9274
rect 7864 9222 7916 9274
rect 12047 9222 12099 9274
rect 12111 9222 12163 9274
rect 12175 9222 12227 9274
rect 12239 9222 12291 9274
rect 12303 9222 12355 9274
rect 16486 9222 16538 9274
rect 16550 9222 16602 9274
rect 16614 9222 16666 9274
rect 16678 9222 16730 9274
rect 16742 9222 16794 9274
rect 5388 8678 5440 8730
rect 5452 8678 5504 8730
rect 5516 8678 5568 8730
rect 5580 8678 5632 8730
rect 5644 8678 5696 8730
rect 9827 8678 9879 8730
rect 9891 8678 9943 8730
rect 9955 8678 10007 8730
rect 10019 8678 10071 8730
rect 10083 8678 10135 8730
rect 14266 8678 14318 8730
rect 14330 8678 14382 8730
rect 14394 8678 14446 8730
rect 14458 8678 14510 8730
rect 14522 8678 14574 8730
rect 18705 8678 18757 8730
rect 18769 8678 18821 8730
rect 18833 8678 18885 8730
rect 18897 8678 18949 8730
rect 18961 8678 19013 8730
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 16948 8508 17000 8560
rect 17132 8440 17184 8492
rect 15936 8372 15988 8424
rect 15752 8347 15804 8356
rect 15752 8313 15761 8347
rect 15761 8313 15795 8347
rect 15795 8313 15804 8347
rect 15752 8304 15804 8313
rect 3169 8134 3221 8186
rect 3233 8134 3285 8186
rect 3297 8134 3349 8186
rect 3361 8134 3413 8186
rect 3425 8134 3477 8186
rect 7608 8134 7660 8186
rect 7672 8134 7724 8186
rect 7736 8134 7788 8186
rect 7800 8134 7852 8186
rect 7864 8134 7916 8186
rect 12047 8134 12099 8186
rect 12111 8134 12163 8186
rect 12175 8134 12227 8186
rect 12239 8134 12291 8186
rect 12303 8134 12355 8186
rect 16486 8134 16538 8186
rect 16550 8134 16602 8186
rect 16614 8134 16666 8186
rect 16678 8134 16730 8186
rect 16742 8134 16794 8186
rect 17040 8032 17092 8084
rect 15936 7964 15988 8016
rect 16396 7964 16448 8016
rect 16948 7896 17000 7948
rect 14924 7692 14976 7744
rect 16764 7871 16816 7880
rect 16764 7837 16773 7871
rect 16773 7837 16807 7871
rect 16807 7837 16816 7871
rect 16764 7828 16816 7837
rect 18420 7939 18472 7948
rect 18420 7905 18429 7939
rect 18429 7905 18463 7939
rect 18463 7905 18472 7939
rect 18420 7896 18472 7905
rect 16120 7735 16172 7744
rect 16120 7701 16129 7735
rect 16129 7701 16163 7735
rect 16163 7701 16172 7735
rect 16120 7692 16172 7701
rect 17408 7735 17460 7744
rect 17408 7701 17417 7735
rect 17417 7701 17451 7735
rect 17451 7701 17460 7735
rect 17408 7692 17460 7701
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 18144 7692 18196 7744
rect 5388 7590 5440 7642
rect 5452 7590 5504 7642
rect 5516 7590 5568 7642
rect 5580 7590 5632 7642
rect 5644 7590 5696 7642
rect 9827 7590 9879 7642
rect 9891 7590 9943 7642
rect 9955 7590 10007 7642
rect 10019 7590 10071 7642
rect 10083 7590 10135 7642
rect 14266 7590 14318 7642
rect 14330 7590 14382 7642
rect 14394 7590 14446 7642
rect 14458 7590 14510 7642
rect 14522 7590 14574 7642
rect 18705 7590 18757 7642
rect 18769 7590 18821 7642
rect 18833 7590 18885 7642
rect 18897 7590 18949 7642
rect 18961 7590 19013 7642
rect 14924 7531 14976 7540
rect 14924 7497 14933 7531
rect 14933 7497 14967 7531
rect 14967 7497 14976 7531
rect 14924 7488 14976 7497
rect 16120 7488 16172 7540
rect 18420 7488 18472 7540
rect 17592 7352 17644 7404
rect 16120 7148 16172 7200
rect 3169 7046 3221 7098
rect 3233 7046 3285 7098
rect 3297 7046 3349 7098
rect 3361 7046 3413 7098
rect 3425 7046 3477 7098
rect 7608 7046 7660 7098
rect 7672 7046 7724 7098
rect 7736 7046 7788 7098
rect 7800 7046 7852 7098
rect 7864 7046 7916 7098
rect 12047 7046 12099 7098
rect 12111 7046 12163 7098
rect 12175 7046 12227 7098
rect 12239 7046 12291 7098
rect 12303 7046 12355 7098
rect 16486 7046 16538 7098
rect 16550 7046 16602 7098
rect 16614 7046 16666 7098
rect 16678 7046 16730 7098
rect 16742 7046 16794 7098
rect 16396 6944 16448 6996
rect 15752 6808 15804 6860
rect 16948 6876 17000 6928
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 17592 6987 17644 6996
rect 17592 6953 17601 6987
rect 17601 6953 17635 6987
rect 17635 6953 17644 6987
rect 17592 6944 17644 6953
rect 17684 6876 17736 6928
rect 18144 6851 18196 6860
rect 18144 6817 18153 6851
rect 18153 6817 18187 6851
rect 18187 6817 18196 6851
rect 18144 6808 18196 6817
rect 16672 6783 16724 6792
rect 16672 6749 16681 6783
rect 16681 6749 16715 6783
rect 16715 6749 16724 6783
rect 16672 6740 16724 6749
rect 16028 6672 16080 6724
rect 17132 6740 17184 6792
rect 16856 6604 16908 6656
rect 5388 6502 5440 6554
rect 5452 6502 5504 6554
rect 5516 6502 5568 6554
rect 5580 6502 5632 6554
rect 5644 6502 5696 6554
rect 9827 6502 9879 6554
rect 9891 6502 9943 6554
rect 9955 6502 10007 6554
rect 10019 6502 10071 6554
rect 10083 6502 10135 6554
rect 14266 6502 14318 6554
rect 14330 6502 14382 6554
rect 14394 6502 14446 6554
rect 14458 6502 14510 6554
rect 14522 6502 14574 6554
rect 18705 6502 18757 6554
rect 18769 6502 18821 6554
rect 18833 6502 18885 6554
rect 18897 6502 18949 6554
rect 18961 6502 19013 6554
rect 16672 6400 16724 6452
rect 17224 6400 17276 6452
rect 3169 5958 3221 6010
rect 3233 5958 3285 6010
rect 3297 5958 3349 6010
rect 3361 5958 3413 6010
rect 3425 5958 3477 6010
rect 7608 5958 7660 6010
rect 7672 5958 7724 6010
rect 7736 5958 7788 6010
rect 7800 5958 7852 6010
rect 7864 5958 7916 6010
rect 12047 5958 12099 6010
rect 12111 5958 12163 6010
rect 12175 5958 12227 6010
rect 12239 5958 12291 6010
rect 12303 5958 12355 6010
rect 16486 5958 16538 6010
rect 16550 5958 16602 6010
rect 16614 5958 16666 6010
rect 16678 5958 16730 6010
rect 16742 5958 16794 6010
rect 16120 5899 16172 5908
rect 16120 5865 16129 5899
rect 16129 5865 16163 5899
rect 16163 5865 16172 5899
rect 16120 5856 16172 5865
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 17408 5584 17460 5593
rect 5388 5414 5440 5466
rect 5452 5414 5504 5466
rect 5516 5414 5568 5466
rect 5580 5414 5632 5466
rect 5644 5414 5696 5466
rect 9827 5414 9879 5466
rect 9891 5414 9943 5466
rect 9955 5414 10007 5466
rect 10019 5414 10071 5466
rect 10083 5414 10135 5466
rect 14266 5414 14318 5466
rect 14330 5414 14382 5466
rect 14394 5414 14446 5466
rect 14458 5414 14510 5466
rect 14522 5414 14574 5466
rect 18705 5414 18757 5466
rect 18769 5414 18821 5466
rect 18833 5414 18885 5466
rect 18897 5414 18949 5466
rect 18961 5414 19013 5466
rect 16396 5312 16448 5364
rect 17040 5312 17092 5364
rect 16028 5244 16080 5296
rect 16304 5176 16356 5228
rect 16856 5176 16908 5228
rect 17684 5108 17736 5160
rect 15936 5015 15988 5024
rect 15936 4981 15945 5015
rect 15945 4981 15979 5015
rect 15979 4981 15988 5015
rect 15936 4972 15988 4981
rect 17408 4972 17460 5024
rect 3169 4870 3221 4922
rect 3233 4870 3285 4922
rect 3297 4870 3349 4922
rect 3361 4870 3413 4922
rect 3425 4870 3477 4922
rect 7608 4870 7660 4922
rect 7672 4870 7724 4922
rect 7736 4870 7788 4922
rect 7800 4870 7852 4922
rect 7864 4870 7916 4922
rect 12047 4870 12099 4922
rect 12111 4870 12163 4922
rect 12175 4870 12227 4922
rect 12239 4870 12291 4922
rect 12303 4870 12355 4922
rect 16486 4870 16538 4922
rect 16550 4870 16602 4922
rect 16614 4870 16666 4922
rect 16678 4870 16730 4922
rect 16742 4870 16794 4922
rect 16028 4539 16080 4548
rect 16028 4505 16062 4539
rect 16062 4505 16080 4539
rect 16028 4496 16080 4505
rect 17316 4607 17368 4616
rect 17316 4573 17325 4607
rect 17325 4573 17359 4607
rect 17359 4573 17368 4607
rect 17316 4564 17368 4573
rect 17684 4564 17736 4616
rect 16120 4428 16172 4480
rect 17132 4471 17184 4480
rect 17132 4437 17141 4471
rect 17141 4437 17175 4471
rect 17175 4437 17184 4471
rect 17132 4428 17184 4437
rect 5388 4326 5440 4378
rect 5452 4326 5504 4378
rect 5516 4326 5568 4378
rect 5580 4326 5632 4378
rect 5644 4326 5696 4378
rect 9827 4326 9879 4378
rect 9891 4326 9943 4378
rect 9955 4326 10007 4378
rect 10019 4326 10071 4378
rect 10083 4326 10135 4378
rect 14266 4326 14318 4378
rect 14330 4326 14382 4378
rect 14394 4326 14446 4378
rect 14458 4326 14510 4378
rect 14522 4326 14574 4378
rect 18705 4326 18757 4378
rect 18769 4326 18821 4378
rect 18833 4326 18885 4378
rect 18897 4326 18949 4378
rect 18961 4326 19013 4378
rect 16028 4224 16080 4276
rect 15936 4088 15988 4140
rect 16304 4131 16356 4140
rect 16304 4097 16313 4131
rect 16313 4097 16347 4131
rect 16347 4097 16356 4131
rect 16304 4088 16356 4097
rect 16396 4131 16448 4140
rect 16396 4097 16405 4131
rect 16405 4097 16439 4131
rect 16439 4097 16448 4131
rect 16396 4088 16448 4097
rect 17684 4088 17736 4140
rect 18328 4063 18380 4072
rect 18328 4029 18337 4063
rect 18337 4029 18371 4063
rect 18371 4029 18380 4063
rect 18328 4020 18380 4029
rect 3169 3782 3221 3834
rect 3233 3782 3285 3834
rect 3297 3782 3349 3834
rect 3361 3782 3413 3834
rect 3425 3782 3477 3834
rect 7608 3782 7660 3834
rect 7672 3782 7724 3834
rect 7736 3782 7788 3834
rect 7800 3782 7852 3834
rect 7864 3782 7916 3834
rect 12047 3782 12099 3834
rect 12111 3782 12163 3834
rect 12175 3782 12227 3834
rect 12239 3782 12291 3834
rect 12303 3782 12355 3834
rect 16486 3782 16538 3834
rect 16550 3782 16602 3834
rect 16614 3782 16666 3834
rect 16678 3782 16730 3834
rect 16742 3782 16794 3834
rect 17316 3680 17368 3732
rect 16396 3612 16448 3664
rect 17132 3544 17184 3596
rect 4988 3476 5040 3528
rect 16856 3476 16908 3528
rect 17408 3519 17460 3528
rect 17408 3485 17417 3519
rect 17417 3485 17451 3519
rect 17451 3485 17460 3519
rect 17408 3476 17460 3485
rect 18420 3451 18472 3460
rect 18420 3417 18429 3451
rect 18429 3417 18463 3451
rect 18463 3417 18472 3451
rect 18420 3408 18472 3417
rect 16120 3383 16172 3392
rect 16120 3349 16129 3383
rect 16129 3349 16163 3383
rect 16163 3349 16172 3383
rect 16120 3340 16172 3349
rect 16488 3340 16540 3392
rect 5388 3238 5440 3290
rect 5452 3238 5504 3290
rect 5516 3238 5568 3290
rect 5580 3238 5632 3290
rect 5644 3238 5696 3290
rect 9827 3238 9879 3290
rect 9891 3238 9943 3290
rect 9955 3238 10007 3290
rect 10019 3238 10071 3290
rect 10083 3238 10135 3290
rect 14266 3238 14318 3290
rect 14330 3238 14382 3290
rect 14394 3238 14446 3290
rect 14458 3238 14510 3290
rect 14522 3238 14574 3290
rect 18705 3238 18757 3290
rect 18769 3238 18821 3290
rect 18833 3238 18885 3290
rect 18897 3238 18949 3290
rect 18961 3238 19013 3290
rect 17684 3136 17736 3188
rect 16212 3000 16264 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 16488 2864 16540 2916
rect 3169 2694 3221 2746
rect 3233 2694 3285 2746
rect 3297 2694 3349 2746
rect 3361 2694 3413 2746
rect 3425 2694 3477 2746
rect 7608 2694 7660 2746
rect 7672 2694 7724 2746
rect 7736 2694 7788 2746
rect 7800 2694 7852 2746
rect 7864 2694 7916 2746
rect 12047 2694 12099 2746
rect 12111 2694 12163 2746
rect 12175 2694 12227 2746
rect 12239 2694 12291 2746
rect 12303 2694 12355 2746
rect 16486 2694 16538 2746
rect 16550 2694 16602 2746
rect 16614 2694 16666 2746
rect 16678 2694 16730 2746
rect 16742 2694 16794 2746
rect 16212 2592 16264 2644
rect 18420 2592 18472 2644
rect 17684 2456 17736 2508
rect 15016 2431 15068 2440
rect 15016 2397 15025 2431
rect 15025 2397 15059 2431
rect 15059 2397 15068 2431
rect 15016 2388 15068 2397
rect 5388 2150 5440 2202
rect 5452 2150 5504 2202
rect 5516 2150 5568 2202
rect 5580 2150 5632 2202
rect 5644 2150 5696 2202
rect 9827 2150 9879 2202
rect 9891 2150 9943 2202
rect 9955 2150 10007 2202
rect 10019 2150 10071 2202
rect 10083 2150 10135 2202
rect 14266 2150 14318 2202
rect 14330 2150 14382 2202
rect 14394 2150 14446 2202
rect 14458 2150 14510 2202
rect 14522 2150 14574 2202
rect 18705 2150 18757 2202
rect 18769 2150 18821 2202
rect 18833 2150 18885 2202
rect 18897 2150 18949 2202
rect 18961 2150 19013 2202
<< metal2 >>
rect 3169 47356 3477 47365
rect 3169 47354 3175 47356
rect 3231 47354 3255 47356
rect 3311 47354 3335 47356
rect 3391 47354 3415 47356
rect 3471 47354 3477 47356
rect 3231 47302 3233 47354
rect 3413 47302 3415 47354
rect 3169 47300 3175 47302
rect 3231 47300 3255 47302
rect 3311 47300 3335 47302
rect 3391 47300 3415 47302
rect 3471 47300 3477 47302
rect 3169 47291 3477 47300
rect 7608 47356 7916 47365
rect 7608 47354 7614 47356
rect 7670 47354 7694 47356
rect 7750 47354 7774 47356
rect 7830 47354 7854 47356
rect 7910 47354 7916 47356
rect 7670 47302 7672 47354
rect 7852 47302 7854 47354
rect 7608 47300 7614 47302
rect 7670 47300 7694 47302
rect 7750 47300 7774 47302
rect 7830 47300 7854 47302
rect 7910 47300 7916 47302
rect 7608 47291 7916 47300
rect 12047 47356 12355 47365
rect 12047 47354 12053 47356
rect 12109 47354 12133 47356
rect 12189 47354 12213 47356
rect 12269 47354 12293 47356
rect 12349 47354 12355 47356
rect 12109 47302 12111 47354
rect 12291 47302 12293 47354
rect 12047 47300 12053 47302
rect 12109 47300 12133 47302
rect 12189 47300 12213 47302
rect 12269 47300 12293 47302
rect 12349 47300 12355 47302
rect 12047 47291 12355 47300
rect 16486 47356 16794 47365
rect 16486 47354 16492 47356
rect 16548 47354 16572 47356
rect 16628 47354 16652 47356
rect 16708 47354 16732 47356
rect 16788 47354 16794 47356
rect 16548 47302 16550 47354
rect 16730 47302 16732 47354
rect 16486 47300 16492 47302
rect 16548 47300 16572 47302
rect 16628 47300 16652 47302
rect 16708 47300 16732 47302
rect 16788 47300 16794 47302
rect 16486 47291 16794 47300
rect 18512 47252 18564 47258
rect 18512 47194 18564 47200
rect 18524 47161 18552 47194
rect 18510 47152 18566 47161
rect 18510 47087 18566 47096
rect 5388 46812 5696 46821
rect 5388 46810 5394 46812
rect 5450 46810 5474 46812
rect 5530 46810 5554 46812
rect 5610 46810 5634 46812
rect 5690 46810 5696 46812
rect 5450 46758 5452 46810
rect 5632 46758 5634 46810
rect 5388 46756 5394 46758
rect 5450 46756 5474 46758
rect 5530 46756 5554 46758
rect 5610 46756 5634 46758
rect 5690 46756 5696 46758
rect 5388 46747 5696 46756
rect 9827 46812 10135 46821
rect 9827 46810 9833 46812
rect 9889 46810 9913 46812
rect 9969 46810 9993 46812
rect 10049 46810 10073 46812
rect 10129 46810 10135 46812
rect 9889 46758 9891 46810
rect 10071 46758 10073 46810
rect 9827 46756 9833 46758
rect 9889 46756 9913 46758
rect 9969 46756 9993 46758
rect 10049 46756 10073 46758
rect 10129 46756 10135 46758
rect 9827 46747 10135 46756
rect 14266 46812 14574 46821
rect 14266 46810 14272 46812
rect 14328 46810 14352 46812
rect 14408 46810 14432 46812
rect 14488 46810 14512 46812
rect 14568 46810 14574 46812
rect 14328 46758 14330 46810
rect 14510 46758 14512 46810
rect 14266 46756 14272 46758
rect 14328 46756 14352 46758
rect 14408 46756 14432 46758
rect 14488 46756 14512 46758
rect 14568 46756 14574 46758
rect 14266 46747 14574 46756
rect 18705 46812 19013 46821
rect 18705 46810 18711 46812
rect 18767 46810 18791 46812
rect 18847 46810 18871 46812
rect 18927 46810 18951 46812
rect 19007 46810 19013 46812
rect 18767 46758 18769 46810
rect 18949 46758 18951 46810
rect 18705 46756 18711 46758
rect 18767 46756 18791 46758
rect 18847 46756 18871 46758
rect 18927 46756 18951 46758
rect 19007 46756 19013 46758
rect 18705 46747 19013 46756
rect 3169 46268 3477 46277
rect 3169 46266 3175 46268
rect 3231 46266 3255 46268
rect 3311 46266 3335 46268
rect 3391 46266 3415 46268
rect 3471 46266 3477 46268
rect 3231 46214 3233 46266
rect 3413 46214 3415 46266
rect 3169 46212 3175 46214
rect 3231 46212 3255 46214
rect 3311 46212 3335 46214
rect 3391 46212 3415 46214
rect 3471 46212 3477 46214
rect 3169 46203 3477 46212
rect 7608 46268 7916 46277
rect 7608 46266 7614 46268
rect 7670 46266 7694 46268
rect 7750 46266 7774 46268
rect 7830 46266 7854 46268
rect 7910 46266 7916 46268
rect 7670 46214 7672 46266
rect 7852 46214 7854 46266
rect 7608 46212 7614 46214
rect 7670 46212 7694 46214
rect 7750 46212 7774 46214
rect 7830 46212 7854 46214
rect 7910 46212 7916 46214
rect 7608 46203 7916 46212
rect 12047 46268 12355 46277
rect 12047 46266 12053 46268
rect 12109 46266 12133 46268
rect 12189 46266 12213 46268
rect 12269 46266 12293 46268
rect 12349 46266 12355 46268
rect 12109 46214 12111 46266
rect 12291 46214 12293 46266
rect 12047 46212 12053 46214
rect 12109 46212 12133 46214
rect 12189 46212 12213 46214
rect 12269 46212 12293 46214
rect 12349 46212 12355 46214
rect 12047 46203 12355 46212
rect 16486 46268 16794 46277
rect 16486 46266 16492 46268
rect 16548 46266 16572 46268
rect 16628 46266 16652 46268
rect 16708 46266 16732 46268
rect 16788 46266 16794 46268
rect 16548 46214 16550 46266
rect 16730 46214 16732 46266
rect 16486 46212 16492 46214
rect 16548 46212 16572 46214
rect 16628 46212 16652 46214
rect 16708 46212 16732 46214
rect 16788 46212 16794 46214
rect 16486 46203 16794 46212
rect 5388 45724 5696 45733
rect 5388 45722 5394 45724
rect 5450 45722 5474 45724
rect 5530 45722 5554 45724
rect 5610 45722 5634 45724
rect 5690 45722 5696 45724
rect 5450 45670 5452 45722
rect 5632 45670 5634 45722
rect 5388 45668 5394 45670
rect 5450 45668 5474 45670
rect 5530 45668 5554 45670
rect 5610 45668 5634 45670
rect 5690 45668 5696 45670
rect 5388 45659 5696 45668
rect 9827 45724 10135 45733
rect 9827 45722 9833 45724
rect 9889 45722 9913 45724
rect 9969 45722 9993 45724
rect 10049 45722 10073 45724
rect 10129 45722 10135 45724
rect 9889 45670 9891 45722
rect 10071 45670 10073 45722
rect 9827 45668 9833 45670
rect 9889 45668 9913 45670
rect 9969 45668 9993 45670
rect 10049 45668 10073 45670
rect 10129 45668 10135 45670
rect 9827 45659 10135 45668
rect 14266 45724 14574 45733
rect 14266 45722 14272 45724
rect 14328 45722 14352 45724
rect 14408 45722 14432 45724
rect 14488 45722 14512 45724
rect 14568 45722 14574 45724
rect 14328 45670 14330 45722
rect 14510 45670 14512 45722
rect 14266 45668 14272 45670
rect 14328 45668 14352 45670
rect 14408 45668 14432 45670
rect 14488 45668 14512 45670
rect 14568 45668 14574 45670
rect 14266 45659 14574 45668
rect 18705 45724 19013 45733
rect 18705 45722 18711 45724
rect 18767 45722 18791 45724
rect 18847 45722 18871 45724
rect 18927 45722 18951 45724
rect 19007 45722 19013 45724
rect 18767 45670 18769 45722
rect 18949 45670 18951 45722
rect 18705 45668 18711 45670
rect 18767 45668 18791 45670
rect 18847 45668 18871 45670
rect 18927 45668 18951 45670
rect 19007 45668 19013 45670
rect 18705 45659 19013 45668
rect 3169 45180 3477 45189
rect 3169 45178 3175 45180
rect 3231 45178 3255 45180
rect 3311 45178 3335 45180
rect 3391 45178 3415 45180
rect 3471 45178 3477 45180
rect 3231 45126 3233 45178
rect 3413 45126 3415 45178
rect 3169 45124 3175 45126
rect 3231 45124 3255 45126
rect 3311 45124 3335 45126
rect 3391 45124 3415 45126
rect 3471 45124 3477 45126
rect 3169 45115 3477 45124
rect 7608 45180 7916 45189
rect 7608 45178 7614 45180
rect 7670 45178 7694 45180
rect 7750 45178 7774 45180
rect 7830 45178 7854 45180
rect 7910 45178 7916 45180
rect 7670 45126 7672 45178
rect 7852 45126 7854 45178
rect 7608 45124 7614 45126
rect 7670 45124 7694 45126
rect 7750 45124 7774 45126
rect 7830 45124 7854 45126
rect 7910 45124 7916 45126
rect 7608 45115 7916 45124
rect 12047 45180 12355 45189
rect 12047 45178 12053 45180
rect 12109 45178 12133 45180
rect 12189 45178 12213 45180
rect 12269 45178 12293 45180
rect 12349 45178 12355 45180
rect 12109 45126 12111 45178
rect 12291 45126 12293 45178
rect 12047 45124 12053 45126
rect 12109 45124 12133 45126
rect 12189 45124 12213 45126
rect 12269 45124 12293 45126
rect 12349 45124 12355 45126
rect 12047 45115 12355 45124
rect 16486 45180 16794 45189
rect 16486 45178 16492 45180
rect 16548 45178 16572 45180
rect 16628 45178 16652 45180
rect 16708 45178 16732 45180
rect 16788 45178 16794 45180
rect 16548 45126 16550 45178
rect 16730 45126 16732 45178
rect 16486 45124 16492 45126
rect 16548 45124 16572 45126
rect 16628 45124 16652 45126
rect 16708 45124 16732 45126
rect 16788 45124 16794 45126
rect 16486 45115 16794 45124
rect 5388 44636 5696 44645
rect 5388 44634 5394 44636
rect 5450 44634 5474 44636
rect 5530 44634 5554 44636
rect 5610 44634 5634 44636
rect 5690 44634 5696 44636
rect 5450 44582 5452 44634
rect 5632 44582 5634 44634
rect 5388 44580 5394 44582
rect 5450 44580 5474 44582
rect 5530 44580 5554 44582
rect 5610 44580 5634 44582
rect 5690 44580 5696 44582
rect 5388 44571 5696 44580
rect 9827 44636 10135 44645
rect 9827 44634 9833 44636
rect 9889 44634 9913 44636
rect 9969 44634 9993 44636
rect 10049 44634 10073 44636
rect 10129 44634 10135 44636
rect 9889 44582 9891 44634
rect 10071 44582 10073 44634
rect 9827 44580 9833 44582
rect 9889 44580 9913 44582
rect 9969 44580 9993 44582
rect 10049 44580 10073 44582
rect 10129 44580 10135 44582
rect 9827 44571 10135 44580
rect 14266 44636 14574 44645
rect 14266 44634 14272 44636
rect 14328 44634 14352 44636
rect 14408 44634 14432 44636
rect 14488 44634 14512 44636
rect 14568 44634 14574 44636
rect 14328 44582 14330 44634
rect 14510 44582 14512 44634
rect 14266 44580 14272 44582
rect 14328 44580 14352 44582
rect 14408 44580 14432 44582
rect 14488 44580 14512 44582
rect 14568 44580 14574 44582
rect 14266 44571 14574 44580
rect 18705 44636 19013 44645
rect 18705 44634 18711 44636
rect 18767 44634 18791 44636
rect 18847 44634 18871 44636
rect 18927 44634 18951 44636
rect 19007 44634 19013 44636
rect 18767 44582 18769 44634
rect 18949 44582 18951 44634
rect 18705 44580 18711 44582
rect 18767 44580 18791 44582
rect 18847 44580 18871 44582
rect 18927 44580 18951 44582
rect 19007 44580 19013 44582
rect 18705 44571 19013 44580
rect 3169 44092 3477 44101
rect 3169 44090 3175 44092
rect 3231 44090 3255 44092
rect 3311 44090 3335 44092
rect 3391 44090 3415 44092
rect 3471 44090 3477 44092
rect 3231 44038 3233 44090
rect 3413 44038 3415 44090
rect 3169 44036 3175 44038
rect 3231 44036 3255 44038
rect 3311 44036 3335 44038
rect 3391 44036 3415 44038
rect 3471 44036 3477 44038
rect 3169 44027 3477 44036
rect 7608 44092 7916 44101
rect 7608 44090 7614 44092
rect 7670 44090 7694 44092
rect 7750 44090 7774 44092
rect 7830 44090 7854 44092
rect 7910 44090 7916 44092
rect 7670 44038 7672 44090
rect 7852 44038 7854 44090
rect 7608 44036 7614 44038
rect 7670 44036 7694 44038
rect 7750 44036 7774 44038
rect 7830 44036 7854 44038
rect 7910 44036 7916 44038
rect 7608 44027 7916 44036
rect 12047 44092 12355 44101
rect 12047 44090 12053 44092
rect 12109 44090 12133 44092
rect 12189 44090 12213 44092
rect 12269 44090 12293 44092
rect 12349 44090 12355 44092
rect 12109 44038 12111 44090
rect 12291 44038 12293 44090
rect 12047 44036 12053 44038
rect 12109 44036 12133 44038
rect 12189 44036 12213 44038
rect 12269 44036 12293 44038
rect 12349 44036 12355 44038
rect 12047 44027 12355 44036
rect 16486 44092 16794 44101
rect 16486 44090 16492 44092
rect 16548 44090 16572 44092
rect 16628 44090 16652 44092
rect 16708 44090 16732 44092
rect 16788 44090 16794 44092
rect 16548 44038 16550 44090
rect 16730 44038 16732 44090
rect 16486 44036 16492 44038
rect 16548 44036 16572 44038
rect 16628 44036 16652 44038
rect 16708 44036 16732 44038
rect 16788 44036 16794 44038
rect 16486 44027 16794 44036
rect 5388 43548 5696 43557
rect 5388 43546 5394 43548
rect 5450 43546 5474 43548
rect 5530 43546 5554 43548
rect 5610 43546 5634 43548
rect 5690 43546 5696 43548
rect 5450 43494 5452 43546
rect 5632 43494 5634 43546
rect 5388 43492 5394 43494
rect 5450 43492 5474 43494
rect 5530 43492 5554 43494
rect 5610 43492 5634 43494
rect 5690 43492 5696 43494
rect 5388 43483 5696 43492
rect 9827 43548 10135 43557
rect 9827 43546 9833 43548
rect 9889 43546 9913 43548
rect 9969 43546 9993 43548
rect 10049 43546 10073 43548
rect 10129 43546 10135 43548
rect 9889 43494 9891 43546
rect 10071 43494 10073 43546
rect 9827 43492 9833 43494
rect 9889 43492 9913 43494
rect 9969 43492 9993 43494
rect 10049 43492 10073 43494
rect 10129 43492 10135 43494
rect 9827 43483 10135 43492
rect 14266 43548 14574 43557
rect 14266 43546 14272 43548
rect 14328 43546 14352 43548
rect 14408 43546 14432 43548
rect 14488 43546 14512 43548
rect 14568 43546 14574 43548
rect 14328 43494 14330 43546
rect 14510 43494 14512 43546
rect 14266 43492 14272 43494
rect 14328 43492 14352 43494
rect 14408 43492 14432 43494
rect 14488 43492 14512 43494
rect 14568 43492 14574 43494
rect 14266 43483 14574 43492
rect 18705 43548 19013 43557
rect 18705 43546 18711 43548
rect 18767 43546 18791 43548
rect 18847 43546 18871 43548
rect 18927 43546 18951 43548
rect 19007 43546 19013 43548
rect 18767 43494 18769 43546
rect 18949 43494 18951 43546
rect 18705 43492 18711 43494
rect 18767 43492 18791 43494
rect 18847 43492 18871 43494
rect 18927 43492 18951 43494
rect 19007 43492 19013 43494
rect 18705 43483 19013 43492
rect 3169 43004 3477 43013
rect 3169 43002 3175 43004
rect 3231 43002 3255 43004
rect 3311 43002 3335 43004
rect 3391 43002 3415 43004
rect 3471 43002 3477 43004
rect 3231 42950 3233 43002
rect 3413 42950 3415 43002
rect 3169 42948 3175 42950
rect 3231 42948 3255 42950
rect 3311 42948 3335 42950
rect 3391 42948 3415 42950
rect 3471 42948 3477 42950
rect 3169 42939 3477 42948
rect 7608 43004 7916 43013
rect 7608 43002 7614 43004
rect 7670 43002 7694 43004
rect 7750 43002 7774 43004
rect 7830 43002 7854 43004
rect 7910 43002 7916 43004
rect 7670 42950 7672 43002
rect 7852 42950 7854 43002
rect 7608 42948 7614 42950
rect 7670 42948 7694 42950
rect 7750 42948 7774 42950
rect 7830 42948 7854 42950
rect 7910 42948 7916 42950
rect 7608 42939 7916 42948
rect 12047 43004 12355 43013
rect 12047 43002 12053 43004
rect 12109 43002 12133 43004
rect 12189 43002 12213 43004
rect 12269 43002 12293 43004
rect 12349 43002 12355 43004
rect 12109 42950 12111 43002
rect 12291 42950 12293 43002
rect 12047 42948 12053 42950
rect 12109 42948 12133 42950
rect 12189 42948 12213 42950
rect 12269 42948 12293 42950
rect 12349 42948 12355 42950
rect 12047 42939 12355 42948
rect 16486 43004 16794 43013
rect 16486 43002 16492 43004
rect 16548 43002 16572 43004
rect 16628 43002 16652 43004
rect 16708 43002 16732 43004
rect 16788 43002 16794 43004
rect 16548 42950 16550 43002
rect 16730 42950 16732 43002
rect 16486 42948 16492 42950
rect 16548 42948 16572 42950
rect 16628 42948 16652 42950
rect 16708 42948 16732 42950
rect 16788 42948 16794 42950
rect 16486 42939 16794 42948
rect 5388 42460 5696 42469
rect 5388 42458 5394 42460
rect 5450 42458 5474 42460
rect 5530 42458 5554 42460
rect 5610 42458 5634 42460
rect 5690 42458 5696 42460
rect 5450 42406 5452 42458
rect 5632 42406 5634 42458
rect 5388 42404 5394 42406
rect 5450 42404 5474 42406
rect 5530 42404 5554 42406
rect 5610 42404 5634 42406
rect 5690 42404 5696 42406
rect 5388 42395 5696 42404
rect 9827 42460 10135 42469
rect 9827 42458 9833 42460
rect 9889 42458 9913 42460
rect 9969 42458 9993 42460
rect 10049 42458 10073 42460
rect 10129 42458 10135 42460
rect 9889 42406 9891 42458
rect 10071 42406 10073 42458
rect 9827 42404 9833 42406
rect 9889 42404 9913 42406
rect 9969 42404 9993 42406
rect 10049 42404 10073 42406
rect 10129 42404 10135 42406
rect 9827 42395 10135 42404
rect 14266 42460 14574 42469
rect 14266 42458 14272 42460
rect 14328 42458 14352 42460
rect 14408 42458 14432 42460
rect 14488 42458 14512 42460
rect 14568 42458 14574 42460
rect 14328 42406 14330 42458
rect 14510 42406 14512 42458
rect 14266 42404 14272 42406
rect 14328 42404 14352 42406
rect 14408 42404 14432 42406
rect 14488 42404 14512 42406
rect 14568 42404 14574 42406
rect 14266 42395 14574 42404
rect 18705 42460 19013 42469
rect 18705 42458 18711 42460
rect 18767 42458 18791 42460
rect 18847 42458 18871 42460
rect 18927 42458 18951 42460
rect 19007 42458 19013 42460
rect 18767 42406 18769 42458
rect 18949 42406 18951 42458
rect 18705 42404 18711 42406
rect 18767 42404 18791 42406
rect 18847 42404 18871 42406
rect 18927 42404 18951 42406
rect 19007 42404 19013 42406
rect 18705 42395 19013 42404
rect 3169 41916 3477 41925
rect 3169 41914 3175 41916
rect 3231 41914 3255 41916
rect 3311 41914 3335 41916
rect 3391 41914 3415 41916
rect 3471 41914 3477 41916
rect 3231 41862 3233 41914
rect 3413 41862 3415 41914
rect 3169 41860 3175 41862
rect 3231 41860 3255 41862
rect 3311 41860 3335 41862
rect 3391 41860 3415 41862
rect 3471 41860 3477 41862
rect 3169 41851 3477 41860
rect 7608 41916 7916 41925
rect 7608 41914 7614 41916
rect 7670 41914 7694 41916
rect 7750 41914 7774 41916
rect 7830 41914 7854 41916
rect 7910 41914 7916 41916
rect 7670 41862 7672 41914
rect 7852 41862 7854 41914
rect 7608 41860 7614 41862
rect 7670 41860 7694 41862
rect 7750 41860 7774 41862
rect 7830 41860 7854 41862
rect 7910 41860 7916 41862
rect 7608 41851 7916 41860
rect 12047 41916 12355 41925
rect 12047 41914 12053 41916
rect 12109 41914 12133 41916
rect 12189 41914 12213 41916
rect 12269 41914 12293 41916
rect 12349 41914 12355 41916
rect 12109 41862 12111 41914
rect 12291 41862 12293 41914
rect 12047 41860 12053 41862
rect 12109 41860 12133 41862
rect 12189 41860 12213 41862
rect 12269 41860 12293 41862
rect 12349 41860 12355 41862
rect 12047 41851 12355 41860
rect 16486 41916 16794 41925
rect 16486 41914 16492 41916
rect 16548 41914 16572 41916
rect 16628 41914 16652 41916
rect 16708 41914 16732 41916
rect 16788 41914 16794 41916
rect 16548 41862 16550 41914
rect 16730 41862 16732 41914
rect 16486 41860 16492 41862
rect 16548 41860 16572 41862
rect 16628 41860 16652 41862
rect 16708 41860 16732 41862
rect 16788 41860 16794 41862
rect 16486 41851 16794 41860
rect 5388 41372 5696 41381
rect 5388 41370 5394 41372
rect 5450 41370 5474 41372
rect 5530 41370 5554 41372
rect 5610 41370 5634 41372
rect 5690 41370 5696 41372
rect 5450 41318 5452 41370
rect 5632 41318 5634 41370
rect 5388 41316 5394 41318
rect 5450 41316 5474 41318
rect 5530 41316 5554 41318
rect 5610 41316 5634 41318
rect 5690 41316 5696 41318
rect 5388 41307 5696 41316
rect 9827 41372 10135 41381
rect 9827 41370 9833 41372
rect 9889 41370 9913 41372
rect 9969 41370 9993 41372
rect 10049 41370 10073 41372
rect 10129 41370 10135 41372
rect 9889 41318 9891 41370
rect 10071 41318 10073 41370
rect 9827 41316 9833 41318
rect 9889 41316 9913 41318
rect 9969 41316 9993 41318
rect 10049 41316 10073 41318
rect 10129 41316 10135 41318
rect 9827 41307 10135 41316
rect 14266 41372 14574 41381
rect 14266 41370 14272 41372
rect 14328 41370 14352 41372
rect 14408 41370 14432 41372
rect 14488 41370 14512 41372
rect 14568 41370 14574 41372
rect 14328 41318 14330 41370
rect 14510 41318 14512 41370
rect 14266 41316 14272 41318
rect 14328 41316 14352 41318
rect 14408 41316 14432 41318
rect 14488 41316 14512 41318
rect 14568 41316 14574 41318
rect 14266 41307 14574 41316
rect 18705 41372 19013 41381
rect 18705 41370 18711 41372
rect 18767 41370 18791 41372
rect 18847 41370 18871 41372
rect 18927 41370 18951 41372
rect 19007 41370 19013 41372
rect 18767 41318 18769 41370
rect 18949 41318 18951 41370
rect 18705 41316 18711 41318
rect 18767 41316 18791 41318
rect 18847 41316 18871 41318
rect 18927 41316 18951 41318
rect 19007 41316 19013 41318
rect 18705 41307 19013 41316
rect 18328 41132 18380 41138
rect 18328 41074 18380 41080
rect 18052 41064 18104 41070
rect 18052 41006 18104 41012
rect 3169 40828 3477 40837
rect 3169 40826 3175 40828
rect 3231 40826 3255 40828
rect 3311 40826 3335 40828
rect 3391 40826 3415 40828
rect 3471 40826 3477 40828
rect 3231 40774 3233 40826
rect 3413 40774 3415 40826
rect 3169 40772 3175 40774
rect 3231 40772 3255 40774
rect 3311 40772 3335 40774
rect 3391 40772 3415 40774
rect 3471 40772 3477 40774
rect 3169 40763 3477 40772
rect 7608 40828 7916 40837
rect 7608 40826 7614 40828
rect 7670 40826 7694 40828
rect 7750 40826 7774 40828
rect 7830 40826 7854 40828
rect 7910 40826 7916 40828
rect 7670 40774 7672 40826
rect 7852 40774 7854 40826
rect 7608 40772 7614 40774
rect 7670 40772 7694 40774
rect 7750 40772 7774 40774
rect 7830 40772 7854 40774
rect 7910 40772 7916 40774
rect 7608 40763 7916 40772
rect 12047 40828 12355 40837
rect 12047 40826 12053 40828
rect 12109 40826 12133 40828
rect 12189 40826 12213 40828
rect 12269 40826 12293 40828
rect 12349 40826 12355 40828
rect 12109 40774 12111 40826
rect 12291 40774 12293 40826
rect 12047 40772 12053 40774
rect 12109 40772 12133 40774
rect 12189 40772 12213 40774
rect 12269 40772 12293 40774
rect 12349 40772 12355 40774
rect 12047 40763 12355 40772
rect 16486 40828 16794 40837
rect 16486 40826 16492 40828
rect 16548 40826 16572 40828
rect 16628 40826 16652 40828
rect 16708 40826 16732 40828
rect 16788 40826 16794 40828
rect 16548 40774 16550 40826
rect 16730 40774 16732 40826
rect 16486 40772 16492 40774
rect 16548 40772 16572 40774
rect 16628 40772 16652 40774
rect 16708 40772 16732 40774
rect 16788 40772 16794 40774
rect 16486 40763 16794 40772
rect 18064 40633 18092 41006
rect 18050 40624 18106 40633
rect 18050 40559 18106 40568
rect 18340 40390 18368 41074
rect 18328 40384 18380 40390
rect 18328 40326 18380 40332
rect 5388 40284 5696 40293
rect 5388 40282 5394 40284
rect 5450 40282 5474 40284
rect 5530 40282 5554 40284
rect 5610 40282 5634 40284
rect 5690 40282 5696 40284
rect 5450 40230 5452 40282
rect 5632 40230 5634 40282
rect 5388 40228 5394 40230
rect 5450 40228 5474 40230
rect 5530 40228 5554 40230
rect 5610 40228 5634 40230
rect 5690 40228 5696 40230
rect 5388 40219 5696 40228
rect 9827 40284 10135 40293
rect 9827 40282 9833 40284
rect 9889 40282 9913 40284
rect 9969 40282 9993 40284
rect 10049 40282 10073 40284
rect 10129 40282 10135 40284
rect 9889 40230 9891 40282
rect 10071 40230 10073 40282
rect 9827 40228 9833 40230
rect 9889 40228 9913 40230
rect 9969 40228 9993 40230
rect 10049 40228 10073 40230
rect 10129 40228 10135 40230
rect 9827 40219 10135 40228
rect 14266 40284 14574 40293
rect 14266 40282 14272 40284
rect 14328 40282 14352 40284
rect 14408 40282 14432 40284
rect 14488 40282 14512 40284
rect 14568 40282 14574 40284
rect 14328 40230 14330 40282
rect 14510 40230 14512 40282
rect 14266 40228 14272 40230
rect 14328 40228 14352 40230
rect 14408 40228 14432 40230
rect 14488 40228 14512 40230
rect 14568 40228 14574 40230
rect 14266 40219 14574 40228
rect 3169 39740 3477 39749
rect 3169 39738 3175 39740
rect 3231 39738 3255 39740
rect 3311 39738 3335 39740
rect 3391 39738 3415 39740
rect 3471 39738 3477 39740
rect 3231 39686 3233 39738
rect 3413 39686 3415 39738
rect 3169 39684 3175 39686
rect 3231 39684 3255 39686
rect 3311 39684 3335 39686
rect 3391 39684 3415 39686
rect 3471 39684 3477 39686
rect 3169 39675 3477 39684
rect 7608 39740 7916 39749
rect 7608 39738 7614 39740
rect 7670 39738 7694 39740
rect 7750 39738 7774 39740
rect 7830 39738 7854 39740
rect 7910 39738 7916 39740
rect 7670 39686 7672 39738
rect 7852 39686 7854 39738
rect 7608 39684 7614 39686
rect 7670 39684 7694 39686
rect 7750 39684 7774 39686
rect 7830 39684 7854 39686
rect 7910 39684 7916 39686
rect 7608 39675 7916 39684
rect 12047 39740 12355 39749
rect 12047 39738 12053 39740
rect 12109 39738 12133 39740
rect 12189 39738 12213 39740
rect 12269 39738 12293 39740
rect 12349 39738 12355 39740
rect 12109 39686 12111 39738
rect 12291 39686 12293 39738
rect 12047 39684 12053 39686
rect 12109 39684 12133 39686
rect 12189 39684 12213 39686
rect 12269 39684 12293 39686
rect 12349 39684 12355 39686
rect 12047 39675 12355 39684
rect 16486 39740 16794 39749
rect 16486 39738 16492 39740
rect 16548 39738 16572 39740
rect 16628 39738 16652 39740
rect 16708 39738 16732 39740
rect 16788 39738 16794 39740
rect 16548 39686 16550 39738
rect 16730 39686 16732 39738
rect 16486 39684 16492 39686
rect 16548 39684 16572 39686
rect 16628 39684 16652 39686
rect 16708 39684 16732 39686
rect 16788 39684 16794 39686
rect 16486 39675 16794 39684
rect 5388 39196 5696 39205
rect 5388 39194 5394 39196
rect 5450 39194 5474 39196
rect 5530 39194 5554 39196
rect 5610 39194 5634 39196
rect 5690 39194 5696 39196
rect 5450 39142 5452 39194
rect 5632 39142 5634 39194
rect 5388 39140 5394 39142
rect 5450 39140 5474 39142
rect 5530 39140 5554 39142
rect 5610 39140 5634 39142
rect 5690 39140 5696 39142
rect 5388 39131 5696 39140
rect 9827 39196 10135 39205
rect 9827 39194 9833 39196
rect 9889 39194 9913 39196
rect 9969 39194 9993 39196
rect 10049 39194 10073 39196
rect 10129 39194 10135 39196
rect 9889 39142 9891 39194
rect 10071 39142 10073 39194
rect 9827 39140 9833 39142
rect 9889 39140 9913 39142
rect 9969 39140 9993 39142
rect 10049 39140 10073 39142
rect 10129 39140 10135 39142
rect 9827 39131 10135 39140
rect 14266 39196 14574 39205
rect 14266 39194 14272 39196
rect 14328 39194 14352 39196
rect 14408 39194 14432 39196
rect 14488 39194 14512 39196
rect 14568 39194 14574 39196
rect 14328 39142 14330 39194
rect 14510 39142 14512 39194
rect 14266 39140 14272 39142
rect 14328 39140 14352 39142
rect 14408 39140 14432 39142
rect 14488 39140 14512 39142
rect 14568 39140 14574 39142
rect 14266 39131 14574 39140
rect 3169 38652 3477 38661
rect 3169 38650 3175 38652
rect 3231 38650 3255 38652
rect 3311 38650 3335 38652
rect 3391 38650 3415 38652
rect 3471 38650 3477 38652
rect 3231 38598 3233 38650
rect 3413 38598 3415 38650
rect 3169 38596 3175 38598
rect 3231 38596 3255 38598
rect 3311 38596 3335 38598
rect 3391 38596 3415 38598
rect 3471 38596 3477 38598
rect 3169 38587 3477 38596
rect 7608 38652 7916 38661
rect 7608 38650 7614 38652
rect 7670 38650 7694 38652
rect 7750 38650 7774 38652
rect 7830 38650 7854 38652
rect 7910 38650 7916 38652
rect 7670 38598 7672 38650
rect 7852 38598 7854 38650
rect 7608 38596 7614 38598
rect 7670 38596 7694 38598
rect 7750 38596 7774 38598
rect 7830 38596 7854 38598
rect 7910 38596 7916 38598
rect 7608 38587 7916 38596
rect 12047 38652 12355 38661
rect 12047 38650 12053 38652
rect 12109 38650 12133 38652
rect 12189 38650 12213 38652
rect 12269 38650 12293 38652
rect 12349 38650 12355 38652
rect 12109 38598 12111 38650
rect 12291 38598 12293 38650
rect 12047 38596 12053 38598
rect 12109 38596 12133 38598
rect 12189 38596 12213 38598
rect 12269 38596 12293 38598
rect 12349 38596 12355 38598
rect 12047 38587 12355 38596
rect 16486 38652 16794 38661
rect 16486 38650 16492 38652
rect 16548 38650 16572 38652
rect 16628 38650 16652 38652
rect 16708 38650 16732 38652
rect 16788 38650 16794 38652
rect 16548 38598 16550 38650
rect 16730 38598 16732 38650
rect 16486 38596 16492 38598
rect 16548 38596 16572 38598
rect 16628 38596 16652 38598
rect 16708 38596 16732 38598
rect 16788 38596 16794 38598
rect 16486 38587 16794 38596
rect 5388 38108 5696 38117
rect 5388 38106 5394 38108
rect 5450 38106 5474 38108
rect 5530 38106 5554 38108
rect 5610 38106 5634 38108
rect 5690 38106 5696 38108
rect 5450 38054 5452 38106
rect 5632 38054 5634 38106
rect 5388 38052 5394 38054
rect 5450 38052 5474 38054
rect 5530 38052 5554 38054
rect 5610 38052 5634 38054
rect 5690 38052 5696 38054
rect 5388 38043 5696 38052
rect 9827 38108 10135 38117
rect 9827 38106 9833 38108
rect 9889 38106 9913 38108
rect 9969 38106 9993 38108
rect 10049 38106 10073 38108
rect 10129 38106 10135 38108
rect 9889 38054 9891 38106
rect 10071 38054 10073 38106
rect 9827 38052 9833 38054
rect 9889 38052 9913 38054
rect 9969 38052 9993 38054
rect 10049 38052 10073 38054
rect 10129 38052 10135 38054
rect 9827 38043 10135 38052
rect 14266 38108 14574 38117
rect 14266 38106 14272 38108
rect 14328 38106 14352 38108
rect 14408 38106 14432 38108
rect 14488 38106 14512 38108
rect 14568 38106 14574 38108
rect 14328 38054 14330 38106
rect 14510 38054 14512 38106
rect 14266 38052 14272 38054
rect 14328 38052 14352 38054
rect 14408 38052 14432 38054
rect 14488 38052 14512 38054
rect 14568 38052 14574 38054
rect 14266 38043 14574 38052
rect 3169 37564 3477 37573
rect 3169 37562 3175 37564
rect 3231 37562 3255 37564
rect 3311 37562 3335 37564
rect 3391 37562 3415 37564
rect 3471 37562 3477 37564
rect 3231 37510 3233 37562
rect 3413 37510 3415 37562
rect 3169 37508 3175 37510
rect 3231 37508 3255 37510
rect 3311 37508 3335 37510
rect 3391 37508 3415 37510
rect 3471 37508 3477 37510
rect 3169 37499 3477 37508
rect 7608 37564 7916 37573
rect 7608 37562 7614 37564
rect 7670 37562 7694 37564
rect 7750 37562 7774 37564
rect 7830 37562 7854 37564
rect 7910 37562 7916 37564
rect 7670 37510 7672 37562
rect 7852 37510 7854 37562
rect 7608 37508 7614 37510
rect 7670 37508 7694 37510
rect 7750 37508 7774 37510
rect 7830 37508 7854 37510
rect 7910 37508 7916 37510
rect 7608 37499 7916 37508
rect 12047 37564 12355 37573
rect 12047 37562 12053 37564
rect 12109 37562 12133 37564
rect 12189 37562 12213 37564
rect 12269 37562 12293 37564
rect 12349 37562 12355 37564
rect 12109 37510 12111 37562
rect 12291 37510 12293 37562
rect 12047 37508 12053 37510
rect 12109 37508 12133 37510
rect 12189 37508 12213 37510
rect 12269 37508 12293 37510
rect 12349 37508 12355 37510
rect 12047 37499 12355 37508
rect 16486 37564 16794 37573
rect 16486 37562 16492 37564
rect 16548 37562 16572 37564
rect 16628 37562 16652 37564
rect 16708 37562 16732 37564
rect 16788 37562 16794 37564
rect 16548 37510 16550 37562
rect 16730 37510 16732 37562
rect 16486 37508 16492 37510
rect 16548 37508 16572 37510
rect 16628 37508 16652 37510
rect 16708 37508 16732 37510
rect 16788 37508 16794 37510
rect 16486 37499 16794 37508
rect 5388 37020 5696 37029
rect 5388 37018 5394 37020
rect 5450 37018 5474 37020
rect 5530 37018 5554 37020
rect 5610 37018 5634 37020
rect 5690 37018 5696 37020
rect 5450 36966 5452 37018
rect 5632 36966 5634 37018
rect 5388 36964 5394 36966
rect 5450 36964 5474 36966
rect 5530 36964 5554 36966
rect 5610 36964 5634 36966
rect 5690 36964 5696 36966
rect 5388 36955 5696 36964
rect 9827 37020 10135 37029
rect 9827 37018 9833 37020
rect 9889 37018 9913 37020
rect 9969 37018 9993 37020
rect 10049 37018 10073 37020
rect 10129 37018 10135 37020
rect 9889 36966 9891 37018
rect 10071 36966 10073 37018
rect 9827 36964 9833 36966
rect 9889 36964 9913 36966
rect 9969 36964 9993 36966
rect 10049 36964 10073 36966
rect 10129 36964 10135 36966
rect 9827 36955 10135 36964
rect 14266 37020 14574 37029
rect 14266 37018 14272 37020
rect 14328 37018 14352 37020
rect 14408 37018 14432 37020
rect 14488 37018 14512 37020
rect 14568 37018 14574 37020
rect 14328 36966 14330 37018
rect 14510 36966 14512 37018
rect 14266 36964 14272 36966
rect 14328 36964 14352 36966
rect 14408 36964 14432 36966
rect 14488 36964 14512 36966
rect 14568 36964 14574 36966
rect 14266 36955 14574 36964
rect 3169 36476 3477 36485
rect 3169 36474 3175 36476
rect 3231 36474 3255 36476
rect 3311 36474 3335 36476
rect 3391 36474 3415 36476
rect 3471 36474 3477 36476
rect 3231 36422 3233 36474
rect 3413 36422 3415 36474
rect 3169 36420 3175 36422
rect 3231 36420 3255 36422
rect 3311 36420 3335 36422
rect 3391 36420 3415 36422
rect 3471 36420 3477 36422
rect 3169 36411 3477 36420
rect 7608 36476 7916 36485
rect 7608 36474 7614 36476
rect 7670 36474 7694 36476
rect 7750 36474 7774 36476
rect 7830 36474 7854 36476
rect 7910 36474 7916 36476
rect 7670 36422 7672 36474
rect 7852 36422 7854 36474
rect 7608 36420 7614 36422
rect 7670 36420 7694 36422
rect 7750 36420 7774 36422
rect 7830 36420 7854 36422
rect 7910 36420 7916 36422
rect 7608 36411 7916 36420
rect 12047 36476 12355 36485
rect 12047 36474 12053 36476
rect 12109 36474 12133 36476
rect 12189 36474 12213 36476
rect 12269 36474 12293 36476
rect 12349 36474 12355 36476
rect 12109 36422 12111 36474
rect 12291 36422 12293 36474
rect 12047 36420 12053 36422
rect 12109 36420 12133 36422
rect 12189 36420 12213 36422
rect 12269 36420 12293 36422
rect 12349 36420 12355 36422
rect 12047 36411 12355 36420
rect 16486 36476 16794 36485
rect 16486 36474 16492 36476
rect 16548 36474 16572 36476
rect 16628 36474 16652 36476
rect 16708 36474 16732 36476
rect 16788 36474 16794 36476
rect 16548 36422 16550 36474
rect 16730 36422 16732 36474
rect 16486 36420 16492 36422
rect 16548 36420 16572 36422
rect 16628 36420 16652 36422
rect 16708 36420 16732 36422
rect 16788 36420 16794 36422
rect 16486 36411 16794 36420
rect 5388 35932 5696 35941
rect 5388 35930 5394 35932
rect 5450 35930 5474 35932
rect 5530 35930 5554 35932
rect 5610 35930 5634 35932
rect 5690 35930 5696 35932
rect 5450 35878 5452 35930
rect 5632 35878 5634 35930
rect 5388 35876 5394 35878
rect 5450 35876 5474 35878
rect 5530 35876 5554 35878
rect 5610 35876 5634 35878
rect 5690 35876 5696 35878
rect 5388 35867 5696 35876
rect 9827 35932 10135 35941
rect 9827 35930 9833 35932
rect 9889 35930 9913 35932
rect 9969 35930 9993 35932
rect 10049 35930 10073 35932
rect 10129 35930 10135 35932
rect 9889 35878 9891 35930
rect 10071 35878 10073 35930
rect 9827 35876 9833 35878
rect 9889 35876 9913 35878
rect 9969 35876 9993 35878
rect 10049 35876 10073 35878
rect 10129 35876 10135 35878
rect 9827 35867 10135 35876
rect 14266 35932 14574 35941
rect 14266 35930 14272 35932
rect 14328 35930 14352 35932
rect 14408 35930 14432 35932
rect 14488 35930 14512 35932
rect 14568 35930 14574 35932
rect 14328 35878 14330 35930
rect 14510 35878 14512 35930
rect 14266 35876 14272 35878
rect 14328 35876 14352 35878
rect 14408 35876 14432 35878
rect 14488 35876 14512 35878
rect 14568 35876 14574 35878
rect 14266 35867 14574 35876
rect 3169 35388 3477 35397
rect 3169 35386 3175 35388
rect 3231 35386 3255 35388
rect 3311 35386 3335 35388
rect 3391 35386 3415 35388
rect 3471 35386 3477 35388
rect 3231 35334 3233 35386
rect 3413 35334 3415 35386
rect 3169 35332 3175 35334
rect 3231 35332 3255 35334
rect 3311 35332 3335 35334
rect 3391 35332 3415 35334
rect 3471 35332 3477 35334
rect 3169 35323 3477 35332
rect 7608 35388 7916 35397
rect 7608 35386 7614 35388
rect 7670 35386 7694 35388
rect 7750 35386 7774 35388
rect 7830 35386 7854 35388
rect 7910 35386 7916 35388
rect 7670 35334 7672 35386
rect 7852 35334 7854 35386
rect 7608 35332 7614 35334
rect 7670 35332 7694 35334
rect 7750 35332 7774 35334
rect 7830 35332 7854 35334
rect 7910 35332 7916 35334
rect 7608 35323 7916 35332
rect 12047 35388 12355 35397
rect 12047 35386 12053 35388
rect 12109 35386 12133 35388
rect 12189 35386 12213 35388
rect 12269 35386 12293 35388
rect 12349 35386 12355 35388
rect 12109 35334 12111 35386
rect 12291 35334 12293 35386
rect 12047 35332 12053 35334
rect 12109 35332 12133 35334
rect 12189 35332 12213 35334
rect 12269 35332 12293 35334
rect 12349 35332 12355 35334
rect 12047 35323 12355 35332
rect 16486 35388 16794 35397
rect 16486 35386 16492 35388
rect 16548 35386 16572 35388
rect 16628 35386 16652 35388
rect 16708 35386 16732 35388
rect 16788 35386 16794 35388
rect 16548 35334 16550 35386
rect 16730 35334 16732 35386
rect 16486 35332 16492 35334
rect 16548 35332 16572 35334
rect 16628 35332 16652 35334
rect 16708 35332 16732 35334
rect 16788 35332 16794 35334
rect 16486 35323 16794 35332
rect 5388 34844 5696 34853
rect 5388 34842 5394 34844
rect 5450 34842 5474 34844
rect 5530 34842 5554 34844
rect 5610 34842 5634 34844
rect 5690 34842 5696 34844
rect 5450 34790 5452 34842
rect 5632 34790 5634 34842
rect 5388 34788 5394 34790
rect 5450 34788 5474 34790
rect 5530 34788 5554 34790
rect 5610 34788 5634 34790
rect 5690 34788 5696 34790
rect 5388 34779 5696 34788
rect 9827 34844 10135 34853
rect 9827 34842 9833 34844
rect 9889 34842 9913 34844
rect 9969 34842 9993 34844
rect 10049 34842 10073 34844
rect 10129 34842 10135 34844
rect 9889 34790 9891 34842
rect 10071 34790 10073 34842
rect 9827 34788 9833 34790
rect 9889 34788 9913 34790
rect 9969 34788 9993 34790
rect 10049 34788 10073 34790
rect 10129 34788 10135 34790
rect 9827 34779 10135 34788
rect 14266 34844 14574 34853
rect 14266 34842 14272 34844
rect 14328 34842 14352 34844
rect 14408 34842 14432 34844
rect 14488 34842 14512 34844
rect 14568 34842 14574 34844
rect 14328 34790 14330 34842
rect 14510 34790 14512 34842
rect 14266 34788 14272 34790
rect 14328 34788 14352 34790
rect 14408 34788 14432 34790
rect 14488 34788 14512 34790
rect 14568 34788 14574 34790
rect 14266 34779 14574 34788
rect 3169 34300 3477 34309
rect 3169 34298 3175 34300
rect 3231 34298 3255 34300
rect 3311 34298 3335 34300
rect 3391 34298 3415 34300
rect 3471 34298 3477 34300
rect 3231 34246 3233 34298
rect 3413 34246 3415 34298
rect 3169 34244 3175 34246
rect 3231 34244 3255 34246
rect 3311 34244 3335 34246
rect 3391 34244 3415 34246
rect 3471 34244 3477 34246
rect 3169 34235 3477 34244
rect 7608 34300 7916 34309
rect 7608 34298 7614 34300
rect 7670 34298 7694 34300
rect 7750 34298 7774 34300
rect 7830 34298 7854 34300
rect 7910 34298 7916 34300
rect 7670 34246 7672 34298
rect 7852 34246 7854 34298
rect 7608 34244 7614 34246
rect 7670 34244 7694 34246
rect 7750 34244 7774 34246
rect 7830 34244 7854 34246
rect 7910 34244 7916 34246
rect 7608 34235 7916 34244
rect 12047 34300 12355 34309
rect 12047 34298 12053 34300
rect 12109 34298 12133 34300
rect 12189 34298 12213 34300
rect 12269 34298 12293 34300
rect 12349 34298 12355 34300
rect 12109 34246 12111 34298
rect 12291 34246 12293 34298
rect 12047 34244 12053 34246
rect 12109 34244 12133 34246
rect 12189 34244 12213 34246
rect 12269 34244 12293 34246
rect 12349 34244 12355 34246
rect 12047 34235 12355 34244
rect 16486 34300 16794 34309
rect 16486 34298 16492 34300
rect 16548 34298 16572 34300
rect 16628 34298 16652 34300
rect 16708 34298 16732 34300
rect 16788 34298 16794 34300
rect 16548 34246 16550 34298
rect 16730 34246 16732 34298
rect 16486 34244 16492 34246
rect 16548 34244 16572 34246
rect 16628 34244 16652 34246
rect 16708 34244 16732 34246
rect 16788 34244 16794 34246
rect 16486 34235 16794 34244
rect 5388 33756 5696 33765
rect 5388 33754 5394 33756
rect 5450 33754 5474 33756
rect 5530 33754 5554 33756
rect 5610 33754 5634 33756
rect 5690 33754 5696 33756
rect 5450 33702 5452 33754
rect 5632 33702 5634 33754
rect 5388 33700 5394 33702
rect 5450 33700 5474 33702
rect 5530 33700 5554 33702
rect 5610 33700 5634 33702
rect 5690 33700 5696 33702
rect 5388 33691 5696 33700
rect 9827 33756 10135 33765
rect 9827 33754 9833 33756
rect 9889 33754 9913 33756
rect 9969 33754 9993 33756
rect 10049 33754 10073 33756
rect 10129 33754 10135 33756
rect 9889 33702 9891 33754
rect 10071 33702 10073 33754
rect 9827 33700 9833 33702
rect 9889 33700 9913 33702
rect 9969 33700 9993 33702
rect 10049 33700 10073 33702
rect 10129 33700 10135 33702
rect 9827 33691 10135 33700
rect 14266 33756 14574 33765
rect 14266 33754 14272 33756
rect 14328 33754 14352 33756
rect 14408 33754 14432 33756
rect 14488 33754 14512 33756
rect 14568 33754 14574 33756
rect 14328 33702 14330 33754
rect 14510 33702 14512 33754
rect 14266 33700 14272 33702
rect 14328 33700 14352 33702
rect 14408 33700 14432 33702
rect 14488 33700 14512 33702
rect 14568 33700 14574 33702
rect 14266 33691 14574 33700
rect 3169 33212 3477 33221
rect 3169 33210 3175 33212
rect 3231 33210 3255 33212
rect 3311 33210 3335 33212
rect 3391 33210 3415 33212
rect 3471 33210 3477 33212
rect 3231 33158 3233 33210
rect 3413 33158 3415 33210
rect 3169 33156 3175 33158
rect 3231 33156 3255 33158
rect 3311 33156 3335 33158
rect 3391 33156 3415 33158
rect 3471 33156 3477 33158
rect 3169 33147 3477 33156
rect 7608 33212 7916 33221
rect 7608 33210 7614 33212
rect 7670 33210 7694 33212
rect 7750 33210 7774 33212
rect 7830 33210 7854 33212
rect 7910 33210 7916 33212
rect 7670 33158 7672 33210
rect 7852 33158 7854 33210
rect 7608 33156 7614 33158
rect 7670 33156 7694 33158
rect 7750 33156 7774 33158
rect 7830 33156 7854 33158
rect 7910 33156 7916 33158
rect 7608 33147 7916 33156
rect 12047 33212 12355 33221
rect 12047 33210 12053 33212
rect 12109 33210 12133 33212
rect 12189 33210 12213 33212
rect 12269 33210 12293 33212
rect 12349 33210 12355 33212
rect 12109 33158 12111 33210
rect 12291 33158 12293 33210
rect 12047 33156 12053 33158
rect 12109 33156 12133 33158
rect 12189 33156 12213 33158
rect 12269 33156 12293 33158
rect 12349 33156 12355 33158
rect 12047 33147 12355 33156
rect 16486 33212 16794 33221
rect 16486 33210 16492 33212
rect 16548 33210 16572 33212
rect 16628 33210 16652 33212
rect 16708 33210 16732 33212
rect 16788 33210 16794 33212
rect 16548 33158 16550 33210
rect 16730 33158 16732 33210
rect 16486 33156 16492 33158
rect 16548 33156 16572 33158
rect 16628 33156 16652 33158
rect 16708 33156 16732 33158
rect 16788 33156 16794 33158
rect 16486 33147 16794 33156
rect 5388 32668 5696 32677
rect 5388 32666 5394 32668
rect 5450 32666 5474 32668
rect 5530 32666 5554 32668
rect 5610 32666 5634 32668
rect 5690 32666 5696 32668
rect 5450 32614 5452 32666
rect 5632 32614 5634 32666
rect 5388 32612 5394 32614
rect 5450 32612 5474 32614
rect 5530 32612 5554 32614
rect 5610 32612 5634 32614
rect 5690 32612 5696 32614
rect 5388 32603 5696 32612
rect 9827 32668 10135 32677
rect 9827 32666 9833 32668
rect 9889 32666 9913 32668
rect 9969 32666 9993 32668
rect 10049 32666 10073 32668
rect 10129 32666 10135 32668
rect 9889 32614 9891 32666
rect 10071 32614 10073 32666
rect 9827 32612 9833 32614
rect 9889 32612 9913 32614
rect 9969 32612 9993 32614
rect 10049 32612 10073 32614
rect 10129 32612 10135 32614
rect 9827 32603 10135 32612
rect 14266 32668 14574 32677
rect 14266 32666 14272 32668
rect 14328 32666 14352 32668
rect 14408 32666 14432 32668
rect 14488 32666 14512 32668
rect 14568 32666 14574 32668
rect 14328 32614 14330 32666
rect 14510 32614 14512 32666
rect 14266 32612 14272 32614
rect 14328 32612 14352 32614
rect 14408 32612 14432 32614
rect 14488 32612 14512 32614
rect 14568 32612 14574 32614
rect 14266 32603 14574 32612
rect 3169 32124 3477 32133
rect 3169 32122 3175 32124
rect 3231 32122 3255 32124
rect 3311 32122 3335 32124
rect 3391 32122 3415 32124
rect 3471 32122 3477 32124
rect 3231 32070 3233 32122
rect 3413 32070 3415 32122
rect 3169 32068 3175 32070
rect 3231 32068 3255 32070
rect 3311 32068 3335 32070
rect 3391 32068 3415 32070
rect 3471 32068 3477 32070
rect 3169 32059 3477 32068
rect 7608 32124 7916 32133
rect 7608 32122 7614 32124
rect 7670 32122 7694 32124
rect 7750 32122 7774 32124
rect 7830 32122 7854 32124
rect 7910 32122 7916 32124
rect 7670 32070 7672 32122
rect 7852 32070 7854 32122
rect 7608 32068 7614 32070
rect 7670 32068 7694 32070
rect 7750 32068 7774 32070
rect 7830 32068 7854 32070
rect 7910 32068 7916 32070
rect 7608 32059 7916 32068
rect 12047 32124 12355 32133
rect 12047 32122 12053 32124
rect 12109 32122 12133 32124
rect 12189 32122 12213 32124
rect 12269 32122 12293 32124
rect 12349 32122 12355 32124
rect 12109 32070 12111 32122
rect 12291 32070 12293 32122
rect 12047 32068 12053 32070
rect 12109 32068 12133 32070
rect 12189 32068 12213 32070
rect 12269 32068 12293 32070
rect 12349 32068 12355 32070
rect 12047 32059 12355 32068
rect 16486 32124 16794 32133
rect 16486 32122 16492 32124
rect 16548 32122 16572 32124
rect 16628 32122 16652 32124
rect 16708 32122 16732 32124
rect 16788 32122 16794 32124
rect 16548 32070 16550 32122
rect 16730 32070 16732 32122
rect 16486 32068 16492 32070
rect 16548 32068 16572 32070
rect 16628 32068 16652 32070
rect 16708 32068 16732 32070
rect 16788 32068 16794 32070
rect 16486 32059 16794 32068
rect 5388 31580 5696 31589
rect 5388 31578 5394 31580
rect 5450 31578 5474 31580
rect 5530 31578 5554 31580
rect 5610 31578 5634 31580
rect 5690 31578 5696 31580
rect 5450 31526 5452 31578
rect 5632 31526 5634 31578
rect 5388 31524 5394 31526
rect 5450 31524 5474 31526
rect 5530 31524 5554 31526
rect 5610 31524 5634 31526
rect 5690 31524 5696 31526
rect 5388 31515 5696 31524
rect 9827 31580 10135 31589
rect 9827 31578 9833 31580
rect 9889 31578 9913 31580
rect 9969 31578 9993 31580
rect 10049 31578 10073 31580
rect 10129 31578 10135 31580
rect 9889 31526 9891 31578
rect 10071 31526 10073 31578
rect 9827 31524 9833 31526
rect 9889 31524 9913 31526
rect 9969 31524 9993 31526
rect 10049 31524 10073 31526
rect 10129 31524 10135 31526
rect 9827 31515 10135 31524
rect 14266 31580 14574 31589
rect 14266 31578 14272 31580
rect 14328 31578 14352 31580
rect 14408 31578 14432 31580
rect 14488 31578 14512 31580
rect 14568 31578 14574 31580
rect 14328 31526 14330 31578
rect 14510 31526 14512 31578
rect 14266 31524 14272 31526
rect 14328 31524 14352 31526
rect 14408 31524 14432 31526
rect 14488 31524 14512 31526
rect 14568 31524 14574 31526
rect 14266 31515 14574 31524
rect 3169 31036 3477 31045
rect 3169 31034 3175 31036
rect 3231 31034 3255 31036
rect 3311 31034 3335 31036
rect 3391 31034 3415 31036
rect 3471 31034 3477 31036
rect 3231 30982 3233 31034
rect 3413 30982 3415 31034
rect 3169 30980 3175 30982
rect 3231 30980 3255 30982
rect 3311 30980 3335 30982
rect 3391 30980 3415 30982
rect 3471 30980 3477 30982
rect 3169 30971 3477 30980
rect 7608 31036 7916 31045
rect 7608 31034 7614 31036
rect 7670 31034 7694 31036
rect 7750 31034 7774 31036
rect 7830 31034 7854 31036
rect 7910 31034 7916 31036
rect 7670 30982 7672 31034
rect 7852 30982 7854 31034
rect 7608 30980 7614 30982
rect 7670 30980 7694 30982
rect 7750 30980 7774 30982
rect 7830 30980 7854 30982
rect 7910 30980 7916 30982
rect 7608 30971 7916 30980
rect 12047 31036 12355 31045
rect 12047 31034 12053 31036
rect 12109 31034 12133 31036
rect 12189 31034 12213 31036
rect 12269 31034 12293 31036
rect 12349 31034 12355 31036
rect 12109 30982 12111 31034
rect 12291 30982 12293 31034
rect 12047 30980 12053 30982
rect 12109 30980 12133 30982
rect 12189 30980 12213 30982
rect 12269 30980 12293 30982
rect 12349 30980 12355 30982
rect 12047 30971 12355 30980
rect 16486 31036 16794 31045
rect 16486 31034 16492 31036
rect 16548 31034 16572 31036
rect 16628 31034 16652 31036
rect 16708 31034 16732 31036
rect 16788 31034 16794 31036
rect 16548 30982 16550 31034
rect 16730 30982 16732 31034
rect 16486 30980 16492 30982
rect 16548 30980 16572 30982
rect 16628 30980 16652 30982
rect 16708 30980 16732 30982
rect 16788 30980 16794 30982
rect 16486 30971 16794 30980
rect 5388 30492 5696 30501
rect 5388 30490 5394 30492
rect 5450 30490 5474 30492
rect 5530 30490 5554 30492
rect 5610 30490 5634 30492
rect 5690 30490 5696 30492
rect 5450 30438 5452 30490
rect 5632 30438 5634 30490
rect 5388 30436 5394 30438
rect 5450 30436 5474 30438
rect 5530 30436 5554 30438
rect 5610 30436 5634 30438
rect 5690 30436 5696 30438
rect 5388 30427 5696 30436
rect 9827 30492 10135 30501
rect 9827 30490 9833 30492
rect 9889 30490 9913 30492
rect 9969 30490 9993 30492
rect 10049 30490 10073 30492
rect 10129 30490 10135 30492
rect 9889 30438 9891 30490
rect 10071 30438 10073 30490
rect 9827 30436 9833 30438
rect 9889 30436 9913 30438
rect 9969 30436 9993 30438
rect 10049 30436 10073 30438
rect 10129 30436 10135 30438
rect 9827 30427 10135 30436
rect 14266 30492 14574 30501
rect 14266 30490 14272 30492
rect 14328 30490 14352 30492
rect 14408 30490 14432 30492
rect 14488 30490 14512 30492
rect 14568 30490 14574 30492
rect 14328 30438 14330 30490
rect 14510 30438 14512 30490
rect 14266 30436 14272 30438
rect 14328 30436 14352 30438
rect 14408 30436 14432 30438
rect 14488 30436 14512 30438
rect 14568 30436 14574 30438
rect 14266 30427 14574 30436
rect 3169 29948 3477 29957
rect 3169 29946 3175 29948
rect 3231 29946 3255 29948
rect 3311 29946 3335 29948
rect 3391 29946 3415 29948
rect 3471 29946 3477 29948
rect 3231 29894 3233 29946
rect 3413 29894 3415 29946
rect 3169 29892 3175 29894
rect 3231 29892 3255 29894
rect 3311 29892 3335 29894
rect 3391 29892 3415 29894
rect 3471 29892 3477 29894
rect 3169 29883 3477 29892
rect 7608 29948 7916 29957
rect 7608 29946 7614 29948
rect 7670 29946 7694 29948
rect 7750 29946 7774 29948
rect 7830 29946 7854 29948
rect 7910 29946 7916 29948
rect 7670 29894 7672 29946
rect 7852 29894 7854 29946
rect 7608 29892 7614 29894
rect 7670 29892 7694 29894
rect 7750 29892 7774 29894
rect 7830 29892 7854 29894
rect 7910 29892 7916 29894
rect 7608 29883 7916 29892
rect 12047 29948 12355 29957
rect 12047 29946 12053 29948
rect 12109 29946 12133 29948
rect 12189 29946 12213 29948
rect 12269 29946 12293 29948
rect 12349 29946 12355 29948
rect 12109 29894 12111 29946
rect 12291 29894 12293 29946
rect 12047 29892 12053 29894
rect 12109 29892 12133 29894
rect 12189 29892 12213 29894
rect 12269 29892 12293 29894
rect 12349 29892 12355 29894
rect 12047 29883 12355 29892
rect 16486 29948 16794 29957
rect 16486 29946 16492 29948
rect 16548 29946 16572 29948
rect 16628 29946 16652 29948
rect 16708 29946 16732 29948
rect 16788 29946 16794 29948
rect 16548 29894 16550 29946
rect 16730 29894 16732 29946
rect 16486 29892 16492 29894
rect 16548 29892 16572 29894
rect 16628 29892 16652 29894
rect 16708 29892 16732 29894
rect 16788 29892 16794 29894
rect 16486 29883 16794 29892
rect 5388 29404 5696 29413
rect 5388 29402 5394 29404
rect 5450 29402 5474 29404
rect 5530 29402 5554 29404
rect 5610 29402 5634 29404
rect 5690 29402 5696 29404
rect 5450 29350 5452 29402
rect 5632 29350 5634 29402
rect 5388 29348 5394 29350
rect 5450 29348 5474 29350
rect 5530 29348 5554 29350
rect 5610 29348 5634 29350
rect 5690 29348 5696 29350
rect 5388 29339 5696 29348
rect 9827 29404 10135 29413
rect 9827 29402 9833 29404
rect 9889 29402 9913 29404
rect 9969 29402 9993 29404
rect 10049 29402 10073 29404
rect 10129 29402 10135 29404
rect 9889 29350 9891 29402
rect 10071 29350 10073 29402
rect 9827 29348 9833 29350
rect 9889 29348 9913 29350
rect 9969 29348 9993 29350
rect 10049 29348 10073 29350
rect 10129 29348 10135 29350
rect 9827 29339 10135 29348
rect 14266 29404 14574 29413
rect 14266 29402 14272 29404
rect 14328 29402 14352 29404
rect 14408 29402 14432 29404
rect 14488 29402 14512 29404
rect 14568 29402 14574 29404
rect 14328 29350 14330 29402
rect 14510 29350 14512 29402
rect 14266 29348 14272 29350
rect 14328 29348 14352 29350
rect 14408 29348 14432 29350
rect 14488 29348 14512 29350
rect 14568 29348 14574 29350
rect 14266 29339 14574 29348
rect 3169 28860 3477 28869
rect 3169 28858 3175 28860
rect 3231 28858 3255 28860
rect 3311 28858 3335 28860
rect 3391 28858 3415 28860
rect 3471 28858 3477 28860
rect 3231 28806 3233 28858
rect 3413 28806 3415 28858
rect 3169 28804 3175 28806
rect 3231 28804 3255 28806
rect 3311 28804 3335 28806
rect 3391 28804 3415 28806
rect 3471 28804 3477 28806
rect 3169 28795 3477 28804
rect 7608 28860 7916 28869
rect 7608 28858 7614 28860
rect 7670 28858 7694 28860
rect 7750 28858 7774 28860
rect 7830 28858 7854 28860
rect 7910 28858 7916 28860
rect 7670 28806 7672 28858
rect 7852 28806 7854 28858
rect 7608 28804 7614 28806
rect 7670 28804 7694 28806
rect 7750 28804 7774 28806
rect 7830 28804 7854 28806
rect 7910 28804 7916 28806
rect 7608 28795 7916 28804
rect 12047 28860 12355 28869
rect 12047 28858 12053 28860
rect 12109 28858 12133 28860
rect 12189 28858 12213 28860
rect 12269 28858 12293 28860
rect 12349 28858 12355 28860
rect 12109 28806 12111 28858
rect 12291 28806 12293 28858
rect 12047 28804 12053 28806
rect 12109 28804 12133 28806
rect 12189 28804 12213 28806
rect 12269 28804 12293 28806
rect 12349 28804 12355 28806
rect 12047 28795 12355 28804
rect 16486 28860 16794 28869
rect 16486 28858 16492 28860
rect 16548 28858 16572 28860
rect 16628 28858 16652 28860
rect 16708 28858 16732 28860
rect 16788 28858 16794 28860
rect 16548 28806 16550 28858
rect 16730 28806 16732 28858
rect 16486 28804 16492 28806
rect 16548 28804 16572 28806
rect 16628 28804 16652 28806
rect 16708 28804 16732 28806
rect 16788 28804 16794 28806
rect 16486 28795 16794 28804
rect 17040 28416 17092 28422
rect 17040 28358 17092 28364
rect 5388 28316 5696 28325
rect 5388 28314 5394 28316
rect 5450 28314 5474 28316
rect 5530 28314 5554 28316
rect 5610 28314 5634 28316
rect 5690 28314 5696 28316
rect 5450 28262 5452 28314
rect 5632 28262 5634 28314
rect 5388 28260 5394 28262
rect 5450 28260 5474 28262
rect 5530 28260 5554 28262
rect 5610 28260 5634 28262
rect 5690 28260 5696 28262
rect 5388 28251 5696 28260
rect 9827 28316 10135 28325
rect 9827 28314 9833 28316
rect 9889 28314 9913 28316
rect 9969 28314 9993 28316
rect 10049 28314 10073 28316
rect 10129 28314 10135 28316
rect 9889 28262 9891 28314
rect 10071 28262 10073 28314
rect 9827 28260 9833 28262
rect 9889 28260 9913 28262
rect 9969 28260 9993 28262
rect 10049 28260 10073 28262
rect 10129 28260 10135 28262
rect 9827 28251 10135 28260
rect 14266 28316 14574 28325
rect 14266 28314 14272 28316
rect 14328 28314 14352 28316
rect 14408 28314 14432 28316
rect 14488 28314 14512 28316
rect 14568 28314 14574 28316
rect 14328 28262 14330 28314
rect 14510 28262 14512 28314
rect 14266 28260 14272 28262
rect 14328 28260 14352 28262
rect 14408 28260 14432 28262
rect 14488 28260 14512 28262
rect 14568 28260 14574 28262
rect 14266 28251 14574 28260
rect 3169 27772 3477 27781
rect 3169 27770 3175 27772
rect 3231 27770 3255 27772
rect 3311 27770 3335 27772
rect 3391 27770 3415 27772
rect 3471 27770 3477 27772
rect 3231 27718 3233 27770
rect 3413 27718 3415 27770
rect 3169 27716 3175 27718
rect 3231 27716 3255 27718
rect 3311 27716 3335 27718
rect 3391 27716 3415 27718
rect 3471 27716 3477 27718
rect 3169 27707 3477 27716
rect 7608 27772 7916 27781
rect 7608 27770 7614 27772
rect 7670 27770 7694 27772
rect 7750 27770 7774 27772
rect 7830 27770 7854 27772
rect 7910 27770 7916 27772
rect 7670 27718 7672 27770
rect 7852 27718 7854 27770
rect 7608 27716 7614 27718
rect 7670 27716 7694 27718
rect 7750 27716 7774 27718
rect 7830 27716 7854 27718
rect 7910 27716 7916 27718
rect 7608 27707 7916 27716
rect 12047 27772 12355 27781
rect 12047 27770 12053 27772
rect 12109 27770 12133 27772
rect 12189 27770 12213 27772
rect 12269 27770 12293 27772
rect 12349 27770 12355 27772
rect 12109 27718 12111 27770
rect 12291 27718 12293 27770
rect 12047 27716 12053 27718
rect 12109 27716 12133 27718
rect 12189 27716 12213 27718
rect 12269 27716 12293 27718
rect 12349 27716 12355 27718
rect 12047 27707 12355 27716
rect 16486 27772 16794 27781
rect 16486 27770 16492 27772
rect 16548 27770 16572 27772
rect 16628 27770 16652 27772
rect 16708 27770 16732 27772
rect 16788 27770 16794 27772
rect 16548 27718 16550 27770
rect 16730 27718 16732 27770
rect 16486 27716 16492 27718
rect 16548 27716 16572 27718
rect 16628 27716 16652 27718
rect 16708 27716 16732 27718
rect 16788 27716 16794 27718
rect 16486 27707 16794 27716
rect 5388 27228 5696 27237
rect 5388 27226 5394 27228
rect 5450 27226 5474 27228
rect 5530 27226 5554 27228
rect 5610 27226 5634 27228
rect 5690 27226 5696 27228
rect 5450 27174 5452 27226
rect 5632 27174 5634 27226
rect 5388 27172 5394 27174
rect 5450 27172 5474 27174
rect 5530 27172 5554 27174
rect 5610 27172 5634 27174
rect 5690 27172 5696 27174
rect 5388 27163 5696 27172
rect 9827 27228 10135 27237
rect 9827 27226 9833 27228
rect 9889 27226 9913 27228
rect 9969 27226 9993 27228
rect 10049 27226 10073 27228
rect 10129 27226 10135 27228
rect 9889 27174 9891 27226
rect 10071 27174 10073 27226
rect 9827 27172 9833 27174
rect 9889 27172 9913 27174
rect 9969 27172 9993 27174
rect 10049 27172 10073 27174
rect 10129 27172 10135 27174
rect 9827 27163 10135 27172
rect 14266 27228 14574 27237
rect 14266 27226 14272 27228
rect 14328 27226 14352 27228
rect 14408 27226 14432 27228
rect 14488 27226 14512 27228
rect 14568 27226 14574 27228
rect 14328 27174 14330 27226
rect 14510 27174 14512 27226
rect 14266 27172 14272 27174
rect 14328 27172 14352 27174
rect 14408 27172 14432 27174
rect 14488 27172 14512 27174
rect 14568 27172 14574 27174
rect 14266 27163 14574 27172
rect 3169 26684 3477 26693
rect 3169 26682 3175 26684
rect 3231 26682 3255 26684
rect 3311 26682 3335 26684
rect 3391 26682 3415 26684
rect 3471 26682 3477 26684
rect 3231 26630 3233 26682
rect 3413 26630 3415 26682
rect 3169 26628 3175 26630
rect 3231 26628 3255 26630
rect 3311 26628 3335 26630
rect 3391 26628 3415 26630
rect 3471 26628 3477 26630
rect 3169 26619 3477 26628
rect 7608 26684 7916 26693
rect 7608 26682 7614 26684
rect 7670 26682 7694 26684
rect 7750 26682 7774 26684
rect 7830 26682 7854 26684
rect 7910 26682 7916 26684
rect 7670 26630 7672 26682
rect 7852 26630 7854 26682
rect 7608 26628 7614 26630
rect 7670 26628 7694 26630
rect 7750 26628 7774 26630
rect 7830 26628 7854 26630
rect 7910 26628 7916 26630
rect 7608 26619 7916 26628
rect 12047 26684 12355 26693
rect 12047 26682 12053 26684
rect 12109 26682 12133 26684
rect 12189 26682 12213 26684
rect 12269 26682 12293 26684
rect 12349 26682 12355 26684
rect 12109 26630 12111 26682
rect 12291 26630 12293 26682
rect 12047 26628 12053 26630
rect 12109 26628 12133 26630
rect 12189 26628 12213 26630
rect 12269 26628 12293 26630
rect 12349 26628 12355 26630
rect 12047 26619 12355 26628
rect 16486 26684 16794 26693
rect 16486 26682 16492 26684
rect 16548 26682 16572 26684
rect 16628 26682 16652 26684
rect 16708 26682 16732 26684
rect 16788 26682 16794 26684
rect 16548 26630 16550 26682
rect 16730 26630 16732 26682
rect 16486 26628 16492 26630
rect 16548 26628 16572 26630
rect 16628 26628 16652 26630
rect 16708 26628 16732 26630
rect 16788 26628 16794 26630
rect 16486 26619 16794 26628
rect 5388 26140 5696 26149
rect 5388 26138 5394 26140
rect 5450 26138 5474 26140
rect 5530 26138 5554 26140
rect 5610 26138 5634 26140
rect 5690 26138 5696 26140
rect 5450 26086 5452 26138
rect 5632 26086 5634 26138
rect 5388 26084 5394 26086
rect 5450 26084 5474 26086
rect 5530 26084 5554 26086
rect 5610 26084 5634 26086
rect 5690 26084 5696 26086
rect 5388 26075 5696 26084
rect 9827 26140 10135 26149
rect 9827 26138 9833 26140
rect 9889 26138 9913 26140
rect 9969 26138 9993 26140
rect 10049 26138 10073 26140
rect 10129 26138 10135 26140
rect 9889 26086 9891 26138
rect 10071 26086 10073 26138
rect 9827 26084 9833 26086
rect 9889 26084 9913 26086
rect 9969 26084 9993 26086
rect 10049 26084 10073 26086
rect 10129 26084 10135 26086
rect 9827 26075 10135 26084
rect 14266 26140 14574 26149
rect 14266 26138 14272 26140
rect 14328 26138 14352 26140
rect 14408 26138 14432 26140
rect 14488 26138 14512 26140
rect 14568 26138 14574 26140
rect 14328 26086 14330 26138
rect 14510 26086 14512 26138
rect 14266 26084 14272 26086
rect 14328 26084 14352 26086
rect 14408 26084 14432 26086
rect 14488 26084 14512 26086
rect 14568 26084 14574 26086
rect 14266 26075 14574 26084
rect 3169 25596 3477 25605
rect 3169 25594 3175 25596
rect 3231 25594 3255 25596
rect 3311 25594 3335 25596
rect 3391 25594 3415 25596
rect 3471 25594 3477 25596
rect 3231 25542 3233 25594
rect 3413 25542 3415 25594
rect 3169 25540 3175 25542
rect 3231 25540 3255 25542
rect 3311 25540 3335 25542
rect 3391 25540 3415 25542
rect 3471 25540 3477 25542
rect 3169 25531 3477 25540
rect 7608 25596 7916 25605
rect 7608 25594 7614 25596
rect 7670 25594 7694 25596
rect 7750 25594 7774 25596
rect 7830 25594 7854 25596
rect 7910 25594 7916 25596
rect 7670 25542 7672 25594
rect 7852 25542 7854 25594
rect 7608 25540 7614 25542
rect 7670 25540 7694 25542
rect 7750 25540 7774 25542
rect 7830 25540 7854 25542
rect 7910 25540 7916 25542
rect 7608 25531 7916 25540
rect 12047 25596 12355 25605
rect 12047 25594 12053 25596
rect 12109 25594 12133 25596
rect 12189 25594 12213 25596
rect 12269 25594 12293 25596
rect 12349 25594 12355 25596
rect 12109 25542 12111 25594
rect 12291 25542 12293 25594
rect 12047 25540 12053 25542
rect 12109 25540 12133 25542
rect 12189 25540 12213 25542
rect 12269 25540 12293 25542
rect 12349 25540 12355 25542
rect 12047 25531 12355 25540
rect 16486 25596 16794 25605
rect 16486 25594 16492 25596
rect 16548 25594 16572 25596
rect 16628 25594 16652 25596
rect 16708 25594 16732 25596
rect 16788 25594 16794 25596
rect 16548 25542 16550 25594
rect 16730 25542 16732 25594
rect 16486 25540 16492 25542
rect 16548 25540 16572 25542
rect 16628 25540 16652 25542
rect 16708 25540 16732 25542
rect 16788 25540 16794 25542
rect 16486 25531 16794 25540
rect 5388 25052 5696 25061
rect 5388 25050 5394 25052
rect 5450 25050 5474 25052
rect 5530 25050 5554 25052
rect 5610 25050 5634 25052
rect 5690 25050 5696 25052
rect 5450 24998 5452 25050
rect 5632 24998 5634 25050
rect 5388 24996 5394 24998
rect 5450 24996 5474 24998
rect 5530 24996 5554 24998
rect 5610 24996 5634 24998
rect 5690 24996 5696 24998
rect 5388 24987 5696 24996
rect 9827 25052 10135 25061
rect 9827 25050 9833 25052
rect 9889 25050 9913 25052
rect 9969 25050 9993 25052
rect 10049 25050 10073 25052
rect 10129 25050 10135 25052
rect 9889 24998 9891 25050
rect 10071 24998 10073 25050
rect 9827 24996 9833 24998
rect 9889 24996 9913 24998
rect 9969 24996 9993 24998
rect 10049 24996 10073 24998
rect 10129 24996 10135 24998
rect 9827 24987 10135 24996
rect 14266 25052 14574 25061
rect 14266 25050 14272 25052
rect 14328 25050 14352 25052
rect 14408 25050 14432 25052
rect 14488 25050 14512 25052
rect 14568 25050 14574 25052
rect 14328 24998 14330 25050
rect 14510 24998 14512 25050
rect 14266 24996 14272 24998
rect 14328 24996 14352 24998
rect 14408 24996 14432 24998
rect 14488 24996 14512 24998
rect 14568 24996 14574 24998
rect 14266 24987 14574 24996
rect 3169 24508 3477 24517
rect 3169 24506 3175 24508
rect 3231 24506 3255 24508
rect 3311 24506 3335 24508
rect 3391 24506 3415 24508
rect 3471 24506 3477 24508
rect 3231 24454 3233 24506
rect 3413 24454 3415 24506
rect 3169 24452 3175 24454
rect 3231 24452 3255 24454
rect 3311 24452 3335 24454
rect 3391 24452 3415 24454
rect 3471 24452 3477 24454
rect 3169 24443 3477 24452
rect 7608 24508 7916 24517
rect 7608 24506 7614 24508
rect 7670 24506 7694 24508
rect 7750 24506 7774 24508
rect 7830 24506 7854 24508
rect 7910 24506 7916 24508
rect 7670 24454 7672 24506
rect 7852 24454 7854 24506
rect 7608 24452 7614 24454
rect 7670 24452 7694 24454
rect 7750 24452 7774 24454
rect 7830 24452 7854 24454
rect 7910 24452 7916 24454
rect 7608 24443 7916 24452
rect 12047 24508 12355 24517
rect 12047 24506 12053 24508
rect 12109 24506 12133 24508
rect 12189 24506 12213 24508
rect 12269 24506 12293 24508
rect 12349 24506 12355 24508
rect 12109 24454 12111 24506
rect 12291 24454 12293 24506
rect 12047 24452 12053 24454
rect 12109 24452 12133 24454
rect 12189 24452 12213 24454
rect 12269 24452 12293 24454
rect 12349 24452 12355 24454
rect 12047 24443 12355 24452
rect 16486 24508 16794 24517
rect 16486 24506 16492 24508
rect 16548 24506 16572 24508
rect 16628 24506 16652 24508
rect 16708 24506 16732 24508
rect 16788 24506 16794 24508
rect 16548 24454 16550 24506
rect 16730 24454 16732 24506
rect 16486 24452 16492 24454
rect 16548 24452 16572 24454
rect 16628 24452 16652 24454
rect 16708 24452 16732 24454
rect 16788 24452 16794 24454
rect 16486 24443 16794 24452
rect 5388 23964 5696 23973
rect 5388 23962 5394 23964
rect 5450 23962 5474 23964
rect 5530 23962 5554 23964
rect 5610 23962 5634 23964
rect 5690 23962 5696 23964
rect 5450 23910 5452 23962
rect 5632 23910 5634 23962
rect 5388 23908 5394 23910
rect 5450 23908 5474 23910
rect 5530 23908 5554 23910
rect 5610 23908 5634 23910
rect 5690 23908 5696 23910
rect 5388 23899 5696 23908
rect 9827 23964 10135 23973
rect 9827 23962 9833 23964
rect 9889 23962 9913 23964
rect 9969 23962 9993 23964
rect 10049 23962 10073 23964
rect 10129 23962 10135 23964
rect 9889 23910 9891 23962
rect 10071 23910 10073 23962
rect 9827 23908 9833 23910
rect 9889 23908 9913 23910
rect 9969 23908 9993 23910
rect 10049 23908 10073 23910
rect 10129 23908 10135 23910
rect 9827 23899 10135 23908
rect 14266 23964 14574 23973
rect 14266 23962 14272 23964
rect 14328 23962 14352 23964
rect 14408 23962 14432 23964
rect 14488 23962 14512 23964
rect 14568 23962 14574 23964
rect 14328 23910 14330 23962
rect 14510 23910 14512 23962
rect 14266 23908 14272 23910
rect 14328 23908 14352 23910
rect 14408 23908 14432 23910
rect 14488 23908 14512 23910
rect 14568 23908 14574 23910
rect 14266 23899 14574 23908
rect 3169 23420 3477 23429
rect 3169 23418 3175 23420
rect 3231 23418 3255 23420
rect 3311 23418 3335 23420
rect 3391 23418 3415 23420
rect 3471 23418 3477 23420
rect 3231 23366 3233 23418
rect 3413 23366 3415 23418
rect 3169 23364 3175 23366
rect 3231 23364 3255 23366
rect 3311 23364 3335 23366
rect 3391 23364 3415 23366
rect 3471 23364 3477 23366
rect 3169 23355 3477 23364
rect 7608 23420 7916 23429
rect 7608 23418 7614 23420
rect 7670 23418 7694 23420
rect 7750 23418 7774 23420
rect 7830 23418 7854 23420
rect 7910 23418 7916 23420
rect 7670 23366 7672 23418
rect 7852 23366 7854 23418
rect 7608 23364 7614 23366
rect 7670 23364 7694 23366
rect 7750 23364 7774 23366
rect 7830 23364 7854 23366
rect 7910 23364 7916 23366
rect 7608 23355 7916 23364
rect 12047 23420 12355 23429
rect 12047 23418 12053 23420
rect 12109 23418 12133 23420
rect 12189 23418 12213 23420
rect 12269 23418 12293 23420
rect 12349 23418 12355 23420
rect 12109 23366 12111 23418
rect 12291 23366 12293 23418
rect 12047 23364 12053 23366
rect 12109 23364 12133 23366
rect 12189 23364 12213 23366
rect 12269 23364 12293 23366
rect 12349 23364 12355 23366
rect 12047 23355 12355 23364
rect 16486 23420 16794 23429
rect 16486 23418 16492 23420
rect 16548 23418 16572 23420
rect 16628 23418 16652 23420
rect 16708 23418 16732 23420
rect 16788 23418 16794 23420
rect 16548 23366 16550 23418
rect 16730 23366 16732 23418
rect 16486 23364 16492 23366
rect 16548 23364 16572 23366
rect 16628 23364 16652 23366
rect 16708 23364 16732 23366
rect 16788 23364 16794 23366
rect 16486 23355 16794 23364
rect 5388 22876 5696 22885
rect 5388 22874 5394 22876
rect 5450 22874 5474 22876
rect 5530 22874 5554 22876
rect 5610 22874 5634 22876
rect 5690 22874 5696 22876
rect 5450 22822 5452 22874
rect 5632 22822 5634 22874
rect 5388 22820 5394 22822
rect 5450 22820 5474 22822
rect 5530 22820 5554 22822
rect 5610 22820 5634 22822
rect 5690 22820 5696 22822
rect 5388 22811 5696 22820
rect 9827 22876 10135 22885
rect 9827 22874 9833 22876
rect 9889 22874 9913 22876
rect 9969 22874 9993 22876
rect 10049 22874 10073 22876
rect 10129 22874 10135 22876
rect 9889 22822 9891 22874
rect 10071 22822 10073 22874
rect 9827 22820 9833 22822
rect 9889 22820 9913 22822
rect 9969 22820 9993 22822
rect 10049 22820 10073 22822
rect 10129 22820 10135 22822
rect 9827 22811 10135 22820
rect 14266 22876 14574 22885
rect 14266 22874 14272 22876
rect 14328 22874 14352 22876
rect 14408 22874 14432 22876
rect 14488 22874 14512 22876
rect 14568 22874 14574 22876
rect 14328 22822 14330 22874
rect 14510 22822 14512 22874
rect 14266 22820 14272 22822
rect 14328 22820 14352 22822
rect 14408 22820 14432 22822
rect 14488 22820 14512 22822
rect 14568 22820 14574 22822
rect 14266 22811 14574 22820
rect 3169 22332 3477 22341
rect 3169 22330 3175 22332
rect 3231 22330 3255 22332
rect 3311 22330 3335 22332
rect 3391 22330 3415 22332
rect 3471 22330 3477 22332
rect 3231 22278 3233 22330
rect 3413 22278 3415 22330
rect 3169 22276 3175 22278
rect 3231 22276 3255 22278
rect 3311 22276 3335 22278
rect 3391 22276 3415 22278
rect 3471 22276 3477 22278
rect 3169 22267 3477 22276
rect 7608 22332 7916 22341
rect 7608 22330 7614 22332
rect 7670 22330 7694 22332
rect 7750 22330 7774 22332
rect 7830 22330 7854 22332
rect 7910 22330 7916 22332
rect 7670 22278 7672 22330
rect 7852 22278 7854 22330
rect 7608 22276 7614 22278
rect 7670 22276 7694 22278
rect 7750 22276 7774 22278
rect 7830 22276 7854 22278
rect 7910 22276 7916 22278
rect 7608 22267 7916 22276
rect 12047 22332 12355 22341
rect 12047 22330 12053 22332
rect 12109 22330 12133 22332
rect 12189 22330 12213 22332
rect 12269 22330 12293 22332
rect 12349 22330 12355 22332
rect 12109 22278 12111 22330
rect 12291 22278 12293 22330
rect 12047 22276 12053 22278
rect 12109 22276 12133 22278
rect 12189 22276 12213 22278
rect 12269 22276 12293 22278
rect 12349 22276 12355 22278
rect 12047 22267 12355 22276
rect 16486 22332 16794 22341
rect 16486 22330 16492 22332
rect 16548 22330 16572 22332
rect 16628 22330 16652 22332
rect 16708 22330 16732 22332
rect 16788 22330 16794 22332
rect 16548 22278 16550 22330
rect 16730 22278 16732 22330
rect 16486 22276 16492 22278
rect 16548 22276 16572 22278
rect 16628 22276 16652 22278
rect 16708 22276 16732 22278
rect 16788 22276 16794 22278
rect 16486 22267 16794 22276
rect 5388 21788 5696 21797
rect 5388 21786 5394 21788
rect 5450 21786 5474 21788
rect 5530 21786 5554 21788
rect 5610 21786 5634 21788
rect 5690 21786 5696 21788
rect 5450 21734 5452 21786
rect 5632 21734 5634 21786
rect 5388 21732 5394 21734
rect 5450 21732 5474 21734
rect 5530 21732 5554 21734
rect 5610 21732 5634 21734
rect 5690 21732 5696 21734
rect 5388 21723 5696 21732
rect 9827 21788 10135 21797
rect 9827 21786 9833 21788
rect 9889 21786 9913 21788
rect 9969 21786 9993 21788
rect 10049 21786 10073 21788
rect 10129 21786 10135 21788
rect 9889 21734 9891 21786
rect 10071 21734 10073 21786
rect 9827 21732 9833 21734
rect 9889 21732 9913 21734
rect 9969 21732 9993 21734
rect 10049 21732 10073 21734
rect 10129 21732 10135 21734
rect 9827 21723 10135 21732
rect 14266 21788 14574 21797
rect 14266 21786 14272 21788
rect 14328 21786 14352 21788
rect 14408 21786 14432 21788
rect 14488 21786 14512 21788
rect 14568 21786 14574 21788
rect 14328 21734 14330 21786
rect 14510 21734 14512 21786
rect 14266 21732 14272 21734
rect 14328 21732 14352 21734
rect 14408 21732 14432 21734
rect 14488 21732 14512 21734
rect 14568 21732 14574 21734
rect 14266 21723 14574 21732
rect 3169 21244 3477 21253
rect 3169 21242 3175 21244
rect 3231 21242 3255 21244
rect 3311 21242 3335 21244
rect 3391 21242 3415 21244
rect 3471 21242 3477 21244
rect 3231 21190 3233 21242
rect 3413 21190 3415 21242
rect 3169 21188 3175 21190
rect 3231 21188 3255 21190
rect 3311 21188 3335 21190
rect 3391 21188 3415 21190
rect 3471 21188 3477 21190
rect 3169 21179 3477 21188
rect 7608 21244 7916 21253
rect 7608 21242 7614 21244
rect 7670 21242 7694 21244
rect 7750 21242 7774 21244
rect 7830 21242 7854 21244
rect 7910 21242 7916 21244
rect 7670 21190 7672 21242
rect 7852 21190 7854 21242
rect 7608 21188 7614 21190
rect 7670 21188 7694 21190
rect 7750 21188 7774 21190
rect 7830 21188 7854 21190
rect 7910 21188 7916 21190
rect 7608 21179 7916 21188
rect 12047 21244 12355 21253
rect 12047 21242 12053 21244
rect 12109 21242 12133 21244
rect 12189 21242 12213 21244
rect 12269 21242 12293 21244
rect 12349 21242 12355 21244
rect 12109 21190 12111 21242
rect 12291 21190 12293 21242
rect 12047 21188 12053 21190
rect 12109 21188 12133 21190
rect 12189 21188 12213 21190
rect 12269 21188 12293 21190
rect 12349 21188 12355 21190
rect 12047 21179 12355 21188
rect 16486 21244 16794 21253
rect 16486 21242 16492 21244
rect 16548 21242 16572 21244
rect 16628 21242 16652 21244
rect 16708 21242 16732 21244
rect 16788 21242 16794 21244
rect 16548 21190 16550 21242
rect 16730 21190 16732 21242
rect 16486 21188 16492 21190
rect 16548 21188 16572 21190
rect 16628 21188 16652 21190
rect 16708 21188 16732 21190
rect 16788 21188 16794 21190
rect 16486 21179 16794 21188
rect 5388 20700 5696 20709
rect 5388 20698 5394 20700
rect 5450 20698 5474 20700
rect 5530 20698 5554 20700
rect 5610 20698 5634 20700
rect 5690 20698 5696 20700
rect 5450 20646 5452 20698
rect 5632 20646 5634 20698
rect 5388 20644 5394 20646
rect 5450 20644 5474 20646
rect 5530 20644 5554 20646
rect 5610 20644 5634 20646
rect 5690 20644 5696 20646
rect 5388 20635 5696 20644
rect 9827 20700 10135 20709
rect 9827 20698 9833 20700
rect 9889 20698 9913 20700
rect 9969 20698 9993 20700
rect 10049 20698 10073 20700
rect 10129 20698 10135 20700
rect 9889 20646 9891 20698
rect 10071 20646 10073 20698
rect 9827 20644 9833 20646
rect 9889 20644 9913 20646
rect 9969 20644 9993 20646
rect 10049 20644 10073 20646
rect 10129 20644 10135 20646
rect 9827 20635 10135 20644
rect 14266 20700 14574 20709
rect 14266 20698 14272 20700
rect 14328 20698 14352 20700
rect 14408 20698 14432 20700
rect 14488 20698 14512 20700
rect 14568 20698 14574 20700
rect 14328 20646 14330 20698
rect 14510 20646 14512 20698
rect 14266 20644 14272 20646
rect 14328 20644 14352 20646
rect 14408 20644 14432 20646
rect 14488 20644 14512 20646
rect 14568 20644 14574 20646
rect 14266 20635 14574 20644
rect 3169 20156 3477 20165
rect 3169 20154 3175 20156
rect 3231 20154 3255 20156
rect 3311 20154 3335 20156
rect 3391 20154 3415 20156
rect 3471 20154 3477 20156
rect 3231 20102 3233 20154
rect 3413 20102 3415 20154
rect 3169 20100 3175 20102
rect 3231 20100 3255 20102
rect 3311 20100 3335 20102
rect 3391 20100 3415 20102
rect 3471 20100 3477 20102
rect 3169 20091 3477 20100
rect 7608 20156 7916 20165
rect 7608 20154 7614 20156
rect 7670 20154 7694 20156
rect 7750 20154 7774 20156
rect 7830 20154 7854 20156
rect 7910 20154 7916 20156
rect 7670 20102 7672 20154
rect 7852 20102 7854 20154
rect 7608 20100 7614 20102
rect 7670 20100 7694 20102
rect 7750 20100 7774 20102
rect 7830 20100 7854 20102
rect 7910 20100 7916 20102
rect 7608 20091 7916 20100
rect 12047 20156 12355 20165
rect 12047 20154 12053 20156
rect 12109 20154 12133 20156
rect 12189 20154 12213 20156
rect 12269 20154 12293 20156
rect 12349 20154 12355 20156
rect 12109 20102 12111 20154
rect 12291 20102 12293 20154
rect 12047 20100 12053 20102
rect 12109 20100 12133 20102
rect 12189 20100 12213 20102
rect 12269 20100 12293 20102
rect 12349 20100 12355 20102
rect 12047 20091 12355 20100
rect 16486 20156 16794 20165
rect 16486 20154 16492 20156
rect 16548 20154 16572 20156
rect 16628 20154 16652 20156
rect 16708 20154 16732 20156
rect 16788 20154 16794 20156
rect 16548 20102 16550 20154
rect 16730 20102 16732 20154
rect 16486 20100 16492 20102
rect 16548 20100 16572 20102
rect 16628 20100 16652 20102
rect 16708 20100 16732 20102
rect 16788 20100 16794 20102
rect 16486 20091 16794 20100
rect 5388 19612 5696 19621
rect 5388 19610 5394 19612
rect 5450 19610 5474 19612
rect 5530 19610 5554 19612
rect 5610 19610 5634 19612
rect 5690 19610 5696 19612
rect 5450 19558 5452 19610
rect 5632 19558 5634 19610
rect 5388 19556 5394 19558
rect 5450 19556 5474 19558
rect 5530 19556 5554 19558
rect 5610 19556 5634 19558
rect 5690 19556 5696 19558
rect 5388 19547 5696 19556
rect 9827 19612 10135 19621
rect 9827 19610 9833 19612
rect 9889 19610 9913 19612
rect 9969 19610 9993 19612
rect 10049 19610 10073 19612
rect 10129 19610 10135 19612
rect 9889 19558 9891 19610
rect 10071 19558 10073 19610
rect 9827 19556 9833 19558
rect 9889 19556 9913 19558
rect 9969 19556 9993 19558
rect 10049 19556 10073 19558
rect 10129 19556 10135 19558
rect 9827 19547 10135 19556
rect 14266 19612 14574 19621
rect 14266 19610 14272 19612
rect 14328 19610 14352 19612
rect 14408 19610 14432 19612
rect 14488 19610 14512 19612
rect 14568 19610 14574 19612
rect 14328 19558 14330 19610
rect 14510 19558 14512 19610
rect 14266 19556 14272 19558
rect 14328 19556 14352 19558
rect 14408 19556 14432 19558
rect 14488 19556 14512 19558
rect 14568 19556 14574 19558
rect 14266 19547 14574 19556
rect 3169 19068 3477 19077
rect 3169 19066 3175 19068
rect 3231 19066 3255 19068
rect 3311 19066 3335 19068
rect 3391 19066 3415 19068
rect 3471 19066 3477 19068
rect 3231 19014 3233 19066
rect 3413 19014 3415 19066
rect 3169 19012 3175 19014
rect 3231 19012 3255 19014
rect 3311 19012 3335 19014
rect 3391 19012 3415 19014
rect 3471 19012 3477 19014
rect 3169 19003 3477 19012
rect 7608 19068 7916 19077
rect 7608 19066 7614 19068
rect 7670 19066 7694 19068
rect 7750 19066 7774 19068
rect 7830 19066 7854 19068
rect 7910 19066 7916 19068
rect 7670 19014 7672 19066
rect 7852 19014 7854 19066
rect 7608 19012 7614 19014
rect 7670 19012 7694 19014
rect 7750 19012 7774 19014
rect 7830 19012 7854 19014
rect 7910 19012 7916 19014
rect 7608 19003 7916 19012
rect 12047 19068 12355 19077
rect 12047 19066 12053 19068
rect 12109 19066 12133 19068
rect 12189 19066 12213 19068
rect 12269 19066 12293 19068
rect 12349 19066 12355 19068
rect 12109 19014 12111 19066
rect 12291 19014 12293 19066
rect 12047 19012 12053 19014
rect 12109 19012 12133 19014
rect 12189 19012 12213 19014
rect 12269 19012 12293 19014
rect 12349 19012 12355 19014
rect 12047 19003 12355 19012
rect 16486 19068 16794 19077
rect 16486 19066 16492 19068
rect 16548 19066 16572 19068
rect 16628 19066 16652 19068
rect 16708 19066 16732 19068
rect 16788 19066 16794 19068
rect 16548 19014 16550 19066
rect 16730 19014 16732 19066
rect 16486 19012 16492 19014
rect 16548 19012 16572 19014
rect 16628 19012 16652 19014
rect 16708 19012 16732 19014
rect 16788 19012 16794 19014
rect 16486 19003 16794 19012
rect 5388 18524 5696 18533
rect 5388 18522 5394 18524
rect 5450 18522 5474 18524
rect 5530 18522 5554 18524
rect 5610 18522 5634 18524
rect 5690 18522 5696 18524
rect 5450 18470 5452 18522
rect 5632 18470 5634 18522
rect 5388 18468 5394 18470
rect 5450 18468 5474 18470
rect 5530 18468 5554 18470
rect 5610 18468 5634 18470
rect 5690 18468 5696 18470
rect 5388 18459 5696 18468
rect 9827 18524 10135 18533
rect 9827 18522 9833 18524
rect 9889 18522 9913 18524
rect 9969 18522 9993 18524
rect 10049 18522 10073 18524
rect 10129 18522 10135 18524
rect 9889 18470 9891 18522
rect 10071 18470 10073 18522
rect 9827 18468 9833 18470
rect 9889 18468 9913 18470
rect 9969 18468 9993 18470
rect 10049 18468 10073 18470
rect 10129 18468 10135 18470
rect 9827 18459 10135 18468
rect 14266 18524 14574 18533
rect 14266 18522 14272 18524
rect 14328 18522 14352 18524
rect 14408 18522 14432 18524
rect 14488 18522 14512 18524
rect 14568 18522 14574 18524
rect 14328 18470 14330 18522
rect 14510 18470 14512 18522
rect 14266 18468 14272 18470
rect 14328 18468 14352 18470
rect 14408 18468 14432 18470
rect 14488 18468 14512 18470
rect 14568 18468 14574 18470
rect 14266 18459 14574 18468
rect 3169 17980 3477 17989
rect 3169 17978 3175 17980
rect 3231 17978 3255 17980
rect 3311 17978 3335 17980
rect 3391 17978 3415 17980
rect 3471 17978 3477 17980
rect 3231 17926 3233 17978
rect 3413 17926 3415 17978
rect 3169 17924 3175 17926
rect 3231 17924 3255 17926
rect 3311 17924 3335 17926
rect 3391 17924 3415 17926
rect 3471 17924 3477 17926
rect 3169 17915 3477 17924
rect 7608 17980 7916 17989
rect 7608 17978 7614 17980
rect 7670 17978 7694 17980
rect 7750 17978 7774 17980
rect 7830 17978 7854 17980
rect 7910 17978 7916 17980
rect 7670 17926 7672 17978
rect 7852 17926 7854 17978
rect 7608 17924 7614 17926
rect 7670 17924 7694 17926
rect 7750 17924 7774 17926
rect 7830 17924 7854 17926
rect 7910 17924 7916 17926
rect 7608 17915 7916 17924
rect 12047 17980 12355 17989
rect 12047 17978 12053 17980
rect 12109 17978 12133 17980
rect 12189 17978 12213 17980
rect 12269 17978 12293 17980
rect 12349 17978 12355 17980
rect 12109 17926 12111 17978
rect 12291 17926 12293 17978
rect 12047 17924 12053 17926
rect 12109 17924 12133 17926
rect 12189 17924 12213 17926
rect 12269 17924 12293 17926
rect 12349 17924 12355 17926
rect 12047 17915 12355 17924
rect 16486 17980 16794 17989
rect 16486 17978 16492 17980
rect 16548 17978 16572 17980
rect 16628 17978 16652 17980
rect 16708 17978 16732 17980
rect 16788 17978 16794 17980
rect 16548 17926 16550 17978
rect 16730 17926 16732 17978
rect 16486 17924 16492 17926
rect 16548 17924 16572 17926
rect 16628 17924 16652 17926
rect 16708 17924 16732 17926
rect 16788 17924 16794 17926
rect 16486 17915 16794 17924
rect 5388 17436 5696 17445
rect 5388 17434 5394 17436
rect 5450 17434 5474 17436
rect 5530 17434 5554 17436
rect 5610 17434 5634 17436
rect 5690 17434 5696 17436
rect 5450 17382 5452 17434
rect 5632 17382 5634 17434
rect 5388 17380 5394 17382
rect 5450 17380 5474 17382
rect 5530 17380 5554 17382
rect 5610 17380 5634 17382
rect 5690 17380 5696 17382
rect 5388 17371 5696 17380
rect 9827 17436 10135 17445
rect 9827 17434 9833 17436
rect 9889 17434 9913 17436
rect 9969 17434 9993 17436
rect 10049 17434 10073 17436
rect 10129 17434 10135 17436
rect 9889 17382 9891 17434
rect 10071 17382 10073 17434
rect 9827 17380 9833 17382
rect 9889 17380 9913 17382
rect 9969 17380 9993 17382
rect 10049 17380 10073 17382
rect 10129 17380 10135 17382
rect 9827 17371 10135 17380
rect 14266 17436 14574 17445
rect 14266 17434 14272 17436
rect 14328 17434 14352 17436
rect 14408 17434 14432 17436
rect 14488 17434 14512 17436
rect 14568 17434 14574 17436
rect 14328 17382 14330 17434
rect 14510 17382 14512 17434
rect 14266 17380 14272 17382
rect 14328 17380 14352 17382
rect 14408 17380 14432 17382
rect 14488 17380 14512 17382
rect 14568 17380 14574 17382
rect 14266 17371 14574 17380
rect 3169 16892 3477 16901
rect 3169 16890 3175 16892
rect 3231 16890 3255 16892
rect 3311 16890 3335 16892
rect 3391 16890 3415 16892
rect 3471 16890 3477 16892
rect 3231 16838 3233 16890
rect 3413 16838 3415 16890
rect 3169 16836 3175 16838
rect 3231 16836 3255 16838
rect 3311 16836 3335 16838
rect 3391 16836 3415 16838
rect 3471 16836 3477 16838
rect 3169 16827 3477 16836
rect 7608 16892 7916 16901
rect 7608 16890 7614 16892
rect 7670 16890 7694 16892
rect 7750 16890 7774 16892
rect 7830 16890 7854 16892
rect 7910 16890 7916 16892
rect 7670 16838 7672 16890
rect 7852 16838 7854 16890
rect 7608 16836 7614 16838
rect 7670 16836 7694 16838
rect 7750 16836 7774 16838
rect 7830 16836 7854 16838
rect 7910 16836 7916 16838
rect 7608 16827 7916 16836
rect 12047 16892 12355 16901
rect 12047 16890 12053 16892
rect 12109 16890 12133 16892
rect 12189 16890 12213 16892
rect 12269 16890 12293 16892
rect 12349 16890 12355 16892
rect 12109 16838 12111 16890
rect 12291 16838 12293 16890
rect 12047 16836 12053 16838
rect 12109 16836 12133 16838
rect 12189 16836 12213 16838
rect 12269 16836 12293 16838
rect 12349 16836 12355 16838
rect 12047 16827 12355 16836
rect 16486 16892 16794 16901
rect 16486 16890 16492 16892
rect 16548 16890 16572 16892
rect 16628 16890 16652 16892
rect 16708 16890 16732 16892
rect 16788 16890 16794 16892
rect 16548 16838 16550 16890
rect 16730 16838 16732 16890
rect 16486 16836 16492 16838
rect 16548 16836 16572 16838
rect 16628 16836 16652 16838
rect 16708 16836 16732 16838
rect 16788 16836 16794 16838
rect 16486 16827 16794 16836
rect 5388 16348 5696 16357
rect 5388 16346 5394 16348
rect 5450 16346 5474 16348
rect 5530 16346 5554 16348
rect 5610 16346 5634 16348
rect 5690 16346 5696 16348
rect 5450 16294 5452 16346
rect 5632 16294 5634 16346
rect 5388 16292 5394 16294
rect 5450 16292 5474 16294
rect 5530 16292 5554 16294
rect 5610 16292 5634 16294
rect 5690 16292 5696 16294
rect 5388 16283 5696 16292
rect 9827 16348 10135 16357
rect 9827 16346 9833 16348
rect 9889 16346 9913 16348
rect 9969 16346 9993 16348
rect 10049 16346 10073 16348
rect 10129 16346 10135 16348
rect 9889 16294 9891 16346
rect 10071 16294 10073 16346
rect 9827 16292 9833 16294
rect 9889 16292 9913 16294
rect 9969 16292 9993 16294
rect 10049 16292 10073 16294
rect 10129 16292 10135 16294
rect 9827 16283 10135 16292
rect 14266 16348 14574 16357
rect 14266 16346 14272 16348
rect 14328 16346 14352 16348
rect 14408 16346 14432 16348
rect 14488 16346 14512 16348
rect 14568 16346 14574 16348
rect 14328 16294 14330 16346
rect 14510 16294 14512 16346
rect 14266 16292 14272 16294
rect 14328 16292 14352 16294
rect 14408 16292 14432 16294
rect 14488 16292 14512 16294
rect 14568 16292 14574 16294
rect 14266 16283 14574 16292
rect 3169 15804 3477 15813
rect 3169 15802 3175 15804
rect 3231 15802 3255 15804
rect 3311 15802 3335 15804
rect 3391 15802 3415 15804
rect 3471 15802 3477 15804
rect 3231 15750 3233 15802
rect 3413 15750 3415 15802
rect 3169 15748 3175 15750
rect 3231 15748 3255 15750
rect 3311 15748 3335 15750
rect 3391 15748 3415 15750
rect 3471 15748 3477 15750
rect 3169 15739 3477 15748
rect 7608 15804 7916 15813
rect 7608 15802 7614 15804
rect 7670 15802 7694 15804
rect 7750 15802 7774 15804
rect 7830 15802 7854 15804
rect 7910 15802 7916 15804
rect 7670 15750 7672 15802
rect 7852 15750 7854 15802
rect 7608 15748 7614 15750
rect 7670 15748 7694 15750
rect 7750 15748 7774 15750
rect 7830 15748 7854 15750
rect 7910 15748 7916 15750
rect 7608 15739 7916 15748
rect 12047 15804 12355 15813
rect 12047 15802 12053 15804
rect 12109 15802 12133 15804
rect 12189 15802 12213 15804
rect 12269 15802 12293 15804
rect 12349 15802 12355 15804
rect 12109 15750 12111 15802
rect 12291 15750 12293 15802
rect 12047 15748 12053 15750
rect 12109 15748 12133 15750
rect 12189 15748 12213 15750
rect 12269 15748 12293 15750
rect 12349 15748 12355 15750
rect 12047 15739 12355 15748
rect 16486 15804 16794 15813
rect 16486 15802 16492 15804
rect 16548 15802 16572 15804
rect 16628 15802 16652 15804
rect 16708 15802 16732 15804
rect 16788 15802 16794 15804
rect 16548 15750 16550 15802
rect 16730 15750 16732 15802
rect 16486 15748 16492 15750
rect 16548 15748 16572 15750
rect 16628 15748 16652 15750
rect 16708 15748 16732 15750
rect 16788 15748 16794 15750
rect 16486 15739 16794 15748
rect 5388 15260 5696 15269
rect 5388 15258 5394 15260
rect 5450 15258 5474 15260
rect 5530 15258 5554 15260
rect 5610 15258 5634 15260
rect 5690 15258 5696 15260
rect 5450 15206 5452 15258
rect 5632 15206 5634 15258
rect 5388 15204 5394 15206
rect 5450 15204 5474 15206
rect 5530 15204 5554 15206
rect 5610 15204 5634 15206
rect 5690 15204 5696 15206
rect 5388 15195 5696 15204
rect 9827 15260 10135 15269
rect 9827 15258 9833 15260
rect 9889 15258 9913 15260
rect 9969 15258 9993 15260
rect 10049 15258 10073 15260
rect 10129 15258 10135 15260
rect 9889 15206 9891 15258
rect 10071 15206 10073 15258
rect 9827 15204 9833 15206
rect 9889 15204 9913 15206
rect 9969 15204 9993 15206
rect 10049 15204 10073 15206
rect 10129 15204 10135 15206
rect 9827 15195 10135 15204
rect 14266 15260 14574 15269
rect 14266 15258 14272 15260
rect 14328 15258 14352 15260
rect 14408 15258 14432 15260
rect 14488 15258 14512 15260
rect 14568 15258 14574 15260
rect 14328 15206 14330 15258
rect 14510 15206 14512 15258
rect 14266 15204 14272 15206
rect 14328 15204 14352 15206
rect 14408 15204 14432 15206
rect 14488 15204 14512 15206
rect 14568 15204 14574 15206
rect 14266 15195 14574 15204
rect 3169 14716 3477 14725
rect 3169 14714 3175 14716
rect 3231 14714 3255 14716
rect 3311 14714 3335 14716
rect 3391 14714 3415 14716
rect 3471 14714 3477 14716
rect 3231 14662 3233 14714
rect 3413 14662 3415 14714
rect 3169 14660 3175 14662
rect 3231 14660 3255 14662
rect 3311 14660 3335 14662
rect 3391 14660 3415 14662
rect 3471 14660 3477 14662
rect 3169 14651 3477 14660
rect 7608 14716 7916 14725
rect 7608 14714 7614 14716
rect 7670 14714 7694 14716
rect 7750 14714 7774 14716
rect 7830 14714 7854 14716
rect 7910 14714 7916 14716
rect 7670 14662 7672 14714
rect 7852 14662 7854 14714
rect 7608 14660 7614 14662
rect 7670 14660 7694 14662
rect 7750 14660 7774 14662
rect 7830 14660 7854 14662
rect 7910 14660 7916 14662
rect 7608 14651 7916 14660
rect 12047 14716 12355 14725
rect 12047 14714 12053 14716
rect 12109 14714 12133 14716
rect 12189 14714 12213 14716
rect 12269 14714 12293 14716
rect 12349 14714 12355 14716
rect 12109 14662 12111 14714
rect 12291 14662 12293 14714
rect 12047 14660 12053 14662
rect 12109 14660 12133 14662
rect 12189 14660 12213 14662
rect 12269 14660 12293 14662
rect 12349 14660 12355 14662
rect 12047 14651 12355 14660
rect 16486 14716 16794 14725
rect 16486 14714 16492 14716
rect 16548 14714 16572 14716
rect 16628 14714 16652 14716
rect 16708 14714 16732 14716
rect 16788 14714 16794 14716
rect 16548 14662 16550 14714
rect 16730 14662 16732 14714
rect 16486 14660 16492 14662
rect 16548 14660 16572 14662
rect 16628 14660 16652 14662
rect 16708 14660 16732 14662
rect 16788 14660 16794 14662
rect 16486 14651 16794 14660
rect 5388 14172 5696 14181
rect 5388 14170 5394 14172
rect 5450 14170 5474 14172
rect 5530 14170 5554 14172
rect 5610 14170 5634 14172
rect 5690 14170 5696 14172
rect 5450 14118 5452 14170
rect 5632 14118 5634 14170
rect 5388 14116 5394 14118
rect 5450 14116 5474 14118
rect 5530 14116 5554 14118
rect 5610 14116 5634 14118
rect 5690 14116 5696 14118
rect 5388 14107 5696 14116
rect 9827 14172 10135 14181
rect 9827 14170 9833 14172
rect 9889 14170 9913 14172
rect 9969 14170 9993 14172
rect 10049 14170 10073 14172
rect 10129 14170 10135 14172
rect 9889 14118 9891 14170
rect 10071 14118 10073 14170
rect 9827 14116 9833 14118
rect 9889 14116 9913 14118
rect 9969 14116 9993 14118
rect 10049 14116 10073 14118
rect 10129 14116 10135 14118
rect 9827 14107 10135 14116
rect 14266 14172 14574 14181
rect 14266 14170 14272 14172
rect 14328 14170 14352 14172
rect 14408 14170 14432 14172
rect 14488 14170 14512 14172
rect 14568 14170 14574 14172
rect 14328 14118 14330 14170
rect 14510 14118 14512 14170
rect 14266 14116 14272 14118
rect 14328 14116 14352 14118
rect 14408 14116 14432 14118
rect 14488 14116 14512 14118
rect 14568 14116 14574 14118
rect 14266 14107 14574 14116
rect 3169 13628 3477 13637
rect 3169 13626 3175 13628
rect 3231 13626 3255 13628
rect 3311 13626 3335 13628
rect 3391 13626 3415 13628
rect 3471 13626 3477 13628
rect 3231 13574 3233 13626
rect 3413 13574 3415 13626
rect 3169 13572 3175 13574
rect 3231 13572 3255 13574
rect 3311 13572 3335 13574
rect 3391 13572 3415 13574
rect 3471 13572 3477 13574
rect 3169 13563 3477 13572
rect 7608 13628 7916 13637
rect 7608 13626 7614 13628
rect 7670 13626 7694 13628
rect 7750 13626 7774 13628
rect 7830 13626 7854 13628
rect 7910 13626 7916 13628
rect 7670 13574 7672 13626
rect 7852 13574 7854 13626
rect 7608 13572 7614 13574
rect 7670 13572 7694 13574
rect 7750 13572 7774 13574
rect 7830 13572 7854 13574
rect 7910 13572 7916 13574
rect 7608 13563 7916 13572
rect 12047 13628 12355 13637
rect 12047 13626 12053 13628
rect 12109 13626 12133 13628
rect 12189 13626 12213 13628
rect 12269 13626 12293 13628
rect 12349 13626 12355 13628
rect 12109 13574 12111 13626
rect 12291 13574 12293 13626
rect 12047 13572 12053 13574
rect 12109 13572 12133 13574
rect 12189 13572 12213 13574
rect 12269 13572 12293 13574
rect 12349 13572 12355 13574
rect 12047 13563 12355 13572
rect 16486 13628 16794 13637
rect 16486 13626 16492 13628
rect 16548 13626 16572 13628
rect 16628 13626 16652 13628
rect 16708 13626 16732 13628
rect 16788 13626 16794 13628
rect 16548 13574 16550 13626
rect 16730 13574 16732 13626
rect 16486 13572 16492 13574
rect 16548 13572 16572 13574
rect 16628 13572 16652 13574
rect 16708 13572 16732 13574
rect 16788 13572 16794 13574
rect 16486 13563 16794 13572
rect 5388 13084 5696 13093
rect 5388 13082 5394 13084
rect 5450 13082 5474 13084
rect 5530 13082 5554 13084
rect 5610 13082 5634 13084
rect 5690 13082 5696 13084
rect 5450 13030 5452 13082
rect 5632 13030 5634 13082
rect 5388 13028 5394 13030
rect 5450 13028 5474 13030
rect 5530 13028 5554 13030
rect 5610 13028 5634 13030
rect 5690 13028 5696 13030
rect 5388 13019 5696 13028
rect 9827 13084 10135 13093
rect 9827 13082 9833 13084
rect 9889 13082 9913 13084
rect 9969 13082 9993 13084
rect 10049 13082 10073 13084
rect 10129 13082 10135 13084
rect 9889 13030 9891 13082
rect 10071 13030 10073 13082
rect 9827 13028 9833 13030
rect 9889 13028 9913 13030
rect 9969 13028 9993 13030
rect 10049 13028 10073 13030
rect 10129 13028 10135 13030
rect 9827 13019 10135 13028
rect 14266 13084 14574 13093
rect 14266 13082 14272 13084
rect 14328 13082 14352 13084
rect 14408 13082 14432 13084
rect 14488 13082 14512 13084
rect 14568 13082 14574 13084
rect 14328 13030 14330 13082
rect 14510 13030 14512 13082
rect 14266 13028 14272 13030
rect 14328 13028 14352 13030
rect 14408 13028 14432 13030
rect 14488 13028 14512 13030
rect 14568 13028 14574 13030
rect 14266 13019 14574 13028
rect 3169 12540 3477 12549
rect 3169 12538 3175 12540
rect 3231 12538 3255 12540
rect 3311 12538 3335 12540
rect 3391 12538 3415 12540
rect 3471 12538 3477 12540
rect 3231 12486 3233 12538
rect 3413 12486 3415 12538
rect 3169 12484 3175 12486
rect 3231 12484 3255 12486
rect 3311 12484 3335 12486
rect 3391 12484 3415 12486
rect 3471 12484 3477 12486
rect 3169 12475 3477 12484
rect 7608 12540 7916 12549
rect 7608 12538 7614 12540
rect 7670 12538 7694 12540
rect 7750 12538 7774 12540
rect 7830 12538 7854 12540
rect 7910 12538 7916 12540
rect 7670 12486 7672 12538
rect 7852 12486 7854 12538
rect 7608 12484 7614 12486
rect 7670 12484 7694 12486
rect 7750 12484 7774 12486
rect 7830 12484 7854 12486
rect 7910 12484 7916 12486
rect 7608 12475 7916 12484
rect 12047 12540 12355 12549
rect 12047 12538 12053 12540
rect 12109 12538 12133 12540
rect 12189 12538 12213 12540
rect 12269 12538 12293 12540
rect 12349 12538 12355 12540
rect 12109 12486 12111 12538
rect 12291 12486 12293 12538
rect 12047 12484 12053 12486
rect 12109 12484 12133 12486
rect 12189 12484 12213 12486
rect 12269 12484 12293 12486
rect 12349 12484 12355 12486
rect 12047 12475 12355 12484
rect 16486 12540 16794 12549
rect 16486 12538 16492 12540
rect 16548 12538 16572 12540
rect 16628 12538 16652 12540
rect 16708 12538 16732 12540
rect 16788 12538 16794 12540
rect 16548 12486 16550 12538
rect 16730 12486 16732 12538
rect 16486 12484 16492 12486
rect 16548 12484 16572 12486
rect 16628 12484 16652 12486
rect 16708 12484 16732 12486
rect 16788 12484 16794 12486
rect 16486 12475 16794 12484
rect 5388 11996 5696 12005
rect 5388 11994 5394 11996
rect 5450 11994 5474 11996
rect 5530 11994 5554 11996
rect 5610 11994 5634 11996
rect 5690 11994 5696 11996
rect 5450 11942 5452 11994
rect 5632 11942 5634 11994
rect 5388 11940 5394 11942
rect 5450 11940 5474 11942
rect 5530 11940 5554 11942
rect 5610 11940 5634 11942
rect 5690 11940 5696 11942
rect 5388 11931 5696 11940
rect 9827 11996 10135 12005
rect 9827 11994 9833 11996
rect 9889 11994 9913 11996
rect 9969 11994 9993 11996
rect 10049 11994 10073 11996
rect 10129 11994 10135 11996
rect 9889 11942 9891 11994
rect 10071 11942 10073 11994
rect 9827 11940 9833 11942
rect 9889 11940 9913 11942
rect 9969 11940 9993 11942
rect 10049 11940 10073 11942
rect 10129 11940 10135 11942
rect 9827 11931 10135 11940
rect 14266 11996 14574 12005
rect 14266 11994 14272 11996
rect 14328 11994 14352 11996
rect 14408 11994 14432 11996
rect 14488 11994 14512 11996
rect 14568 11994 14574 11996
rect 14328 11942 14330 11994
rect 14510 11942 14512 11994
rect 14266 11940 14272 11942
rect 14328 11940 14352 11942
rect 14408 11940 14432 11942
rect 14488 11940 14512 11942
rect 14568 11940 14574 11942
rect 14266 11931 14574 11940
rect 3169 11452 3477 11461
rect 3169 11450 3175 11452
rect 3231 11450 3255 11452
rect 3311 11450 3335 11452
rect 3391 11450 3415 11452
rect 3471 11450 3477 11452
rect 3231 11398 3233 11450
rect 3413 11398 3415 11450
rect 3169 11396 3175 11398
rect 3231 11396 3255 11398
rect 3311 11396 3335 11398
rect 3391 11396 3415 11398
rect 3471 11396 3477 11398
rect 3169 11387 3477 11396
rect 7608 11452 7916 11461
rect 7608 11450 7614 11452
rect 7670 11450 7694 11452
rect 7750 11450 7774 11452
rect 7830 11450 7854 11452
rect 7910 11450 7916 11452
rect 7670 11398 7672 11450
rect 7852 11398 7854 11450
rect 7608 11396 7614 11398
rect 7670 11396 7694 11398
rect 7750 11396 7774 11398
rect 7830 11396 7854 11398
rect 7910 11396 7916 11398
rect 7608 11387 7916 11396
rect 12047 11452 12355 11461
rect 12047 11450 12053 11452
rect 12109 11450 12133 11452
rect 12189 11450 12213 11452
rect 12269 11450 12293 11452
rect 12349 11450 12355 11452
rect 12109 11398 12111 11450
rect 12291 11398 12293 11450
rect 12047 11396 12053 11398
rect 12109 11396 12133 11398
rect 12189 11396 12213 11398
rect 12269 11396 12293 11398
rect 12349 11396 12355 11398
rect 12047 11387 12355 11396
rect 16486 11452 16794 11461
rect 16486 11450 16492 11452
rect 16548 11450 16572 11452
rect 16628 11450 16652 11452
rect 16708 11450 16732 11452
rect 16788 11450 16794 11452
rect 16548 11398 16550 11450
rect 16730 11398 16732 11450
rect 16486 11396 16492 11398
rect 16548 11396 16572 11398
rect 16628 11396 16652 11398
rect 16708 11396 16732 11398
rect 16788 11396 16794 11398
rect 16486 11387 16794 11396
rect 5388 10908 5696 10917
rect 5388 10906 5394 10908
rect 5450 10906 5474 10908
rect 5530 10906 5554 10908
rect 5610 10906 5634 10908
rect 5690 10906 5696 10908
rect 5450 10854 5452 10906
rect 5632 10854 5634 10906
rect 5388 10852 5394 10854
rect 5450 10852 5474 10854
rect 5530 10852 5554 10854
rect 5610 10852 5634 10854
rect 5690 10852 5696 10854
rect 5388 10843 5696 10852
rect 9827 10908 10135 10917
rect 9827 10906 9833 10908
rect 9889 10906 9913 10908
rect 9969 10906 9993 10908
rect 10049 10906 10073 10908
rect 10129 10906 10135 10908
rect 9889 10854 9891 10906
rect 10071 10854 10073 10906
rect 9827 10852 9833 10854
rect 9889 10852 9913 10854
rect 9969 10852 9993 10854
rect 10049 10852 10073 10854
rect 10129 10852 10135 10854
rect 9827 10843 10135 10852
rect 14266 10908 14574 10917
rect 14266 10906 14272 10908
rect 14328 10906 14352 10908
rect 14408 10906 14432 10908
rect 14488 10906 14512 10908
rect 14568 10906 14574 10908
rect 14328 10854 14330 10906
rect 14510 10854 14512 10906
rect 14266 10852 14272 10854
rect 14328 10852 14352 10854
rect 14408 10852 14432 10854
rect 14488 10852 14512 10854
rect 14568 10852 14574 10854
rect 14266 10843 14574 10852
rect 3169 10364 3477 10373
rect 3169 10362 3175 10364
rect 3231 10362 3255 10364
rect 3311 10362 3335 10364
rect 3391 10362 3415 10364
rect 3471 10362 3477 10364
rect 3231 10310 3233 10362
rect 3413 10310 3415 10362
rect 3169 10308 3175 10310
rect 3231 10308 3255 10310
rect 3311 10308 3335 10310
rect 3391 10308 3415 10310
rect 3471 10308 3477 10310
rect 3169 10299 3477 10308
rect 7608 10364 7916 10373
rect 7608 10362 7614 10364
rect 7670 10362 7694 10364
rect 7750 10362 7774 10364
rect 7830 10362 7854 10364
rect 7910 10362 7916 10364
rect 7670 10310 7672 10362
rect 7852 10310 7854 10362
rect 7608 10308 7614 10310
rect 7670 10308 7694 10310
rect 7750 10308 7774 10310
rect 7830 10308 7854 10310
rect 7910 10308 7916 10310
rect 7608 10299 7916 10308
rect 12047 10364 12355 10373
rect 12047 10362 12053 10364
rect 12109 10362 12133 10364
rect 12189 10362 12213 10364
rect 12269 10362 12293 10364
rect 12349 10362 12355 10364
rect 12109 10310 12111 10362
rect 12291 10310 12293 10362
rect 12047 10308 12053 10310
rect 12109 10308 12133 10310
rect 12189 10308 12213 10310
rect 12269 10308 12293 10310
rect 12349 10308 12355 10310
rect 12047 10299 12355 10308
rect 16486 10364 16794 10373
rect 16486 10362 16492 10364
rect 16548 10362 16572 10364
rect 16628 10362 16652 10364
rect 16708 10362 16732 10364
rect 16788 10362 16794 10364
rect 16548 10310 16550 10362
rect 16730 10310 16732 10362
rect 16486 10308 16492 10310
rect 16548 10308 16572 10310
rect 16628 10308 16652 10310
rect 16708 10308 16732 10310
rect 16788 10308 16794 10310
rect 16486 10299 16794 10308
rect 5388 9820 5696 9829
rect 5388 9818 5394 9820
rect 5450 9818 5474 9820
rect 5530 9818 5554 9820
rect 5610 9818 5634 9820
rect 5690 9818 5696 9820
rect 5450 9766 5452 9818
rect 5632 9766 5634 9818
rect 5388 9764 5394 9766
rect 5450 9764 5474 9766
rect 5530 9764 5554 9766
rect 5610 9764 5634 9766
rect 5690 9764 5696 9766
rect 5388 9755 5696 9764
rect 9827 9820 10135 9829
rect 9827 9818 9833 9820
rect 9889 9818 9913 9820
rect 9969 9818 9993 9820
rect 10049 9818 10073 9820
rect 10129 9818 10135 9820
rect 9889 9766 9891 9818
rect 10071 9766 10073 9818
rect 9827 9764 9833 9766
rect 9889 9764 9913 9766
rect 9969 9764 9993 9766
rect 10049 9764 10073 9766
rect 10129 9764 10135 9766
rect 9827 9755 10135 9764
rect 14266 9820 14574 9829
rect 14266 9818 14272 9820
rect 14328 9818 14352 9820
rect 14408 9818 14432 9820
rect 14488 9818 14512 9820
rect 14568 9818 14574 9820
rect 14328 9766 14330 9818
rect 14510 9766 14512 9818
rect 14266 9764 14272 9766
rect 14328 9764 14352 9766
rect 14408 9764 14432 9766
rect 14488 9764 14512 9766
rect 14568 9764 14574 9766
rect 14266 9755 14574 9764
rect 3169 9276 3477 9285
rect 3169 9274 3175 9276
rect 3231 9274 3255 9276
rect 3311 9274 3335 9276
rect 3391 9274 3415 9276
rect 3471 9274 3477 9276
rect 3231 9222 3233 9274
rect 3413 9222 3415 9274
rect 3169 9220 3175 9222
rect 3231 9220 3255 9222
rect 3311 9220 3335 9222
rect 3391 9220 3415 9222
rect 3471 9220 3477 9222
rect 3169 9211 3477 9220
rect 7608 9276 7916 9285
rect 7608 9274 7614 9276
rect 7670 9274 7694 9276
rect 7750 9274 7774 9276
rect 7830 9274 7854 9276
rect 7910 9274 7916 9276
rect 7670 9222 7672 9274
rect 7852 9222 7854 9274
rect 7608 9220 7614 9222
rect 7670 9220 7694 9222
rect 7750 9220 7774 9222
rect 7830 9220 7854 9222
rect 7910 9220 7916 9222
rect 7608 9211 7916 9220
rect 12047 9276 12355 9285
rect 12047 9274 12053 9276
rect 12109 9274 12133 9276
rect 12189 9274 12213 9276
rect 12269 9274 12293 9276
rect 12349 9274 12355 9276
rect 12109 9222 12111 9274
rect 12291 9222 12293 9274
rect 12047 9220 12053 9222
rect 12109 9220 12133 9222
rect 12189 9220 12213 9222
rect 12269 9220 12293 9222
rect 12349 9220 12355 9222
rect 12047 9211 12355 9220
rect 16486 9276 16794 9285
rect 16486 9274 16492 9276
rect 16548 9274 16572 9276
rect 16628 9274 16652 9276
rect 16708 9274 16732 9276
rect 16788 9274 16794 9276
rect 16548 9222 16550 9274
rect 16730 9222 16732 9274
rect 16486 9220 16492 9222
rect 16548 9220 16572 9222
rect 16628 9220 16652 9222
rect 16708 9220 16732 9222
rect 16788 9220 16794 9222
rect 16486 9211 16794 9220
rect 5388 8732 5696 8741
rect 5388 8730 5394 8732
rect 5450 8730 5474 8732
rect 5530 8730 5554 8732
rect 5610 8730 5634 8732
rect 5690 8730 5696 8732
rect 5450 8678 5452 8730
rect 5632 8678 5634 8730
rect 5388 8676 5394 8678
rect 5450 8676 5474 8678
rect 5530 8676 5554 8678
rect 5610 8676 5634 8678
rect 5690 8676 5696 8678
rect 5388 8667 5696 8676
rect 9827 8732 10135 8741
rect 9827 8730 9833 8732
rect 9889 8730 9913 8732
rect 9969 8730 9993 8732
rect 10049 8730 10073 8732
rect 10129 8730 10135 8732
rect 9889 8678 9891 8730
rect 10071 8678 10073 8730
rect 9827 8676 9833 8678
rect 9889 8676 9913 8678
rect 9969 8676 9993 8678
rect 10049 8676 10073 8678
rect 10129 8676 10135 8678
rect 9827 8667 10135 8676
rect 14266 8732 14574 8741
rect 14266 8730 14272 8732
rect 14328 8730 14352 8732
rect 14408 8730 14432 8732
rect 14488 8730 14512 8732
rect 14568 8730 14574 8732
rect 14328 8678 14330 8730
rect 14510 8678 14512 8730
rect 14266 8676 14272 8678
rect 14328 8676 14352 8678
rect 14408 8676 14432 8678
rect 14488 8676 14512 8678
rect 14568 8676 14574 8678
rect 14266 8667 14574 8676
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 15936 8424 15988 8430
rect 15936 8366 15988 8372
rect 15752 8356 15804 8362
rect 15752 8298 15804 8304
rect 3169 8188 3477 8197
rect 3169 8186 3175 8188
rect 3231 8186 3255 8188
rect 3311 8186 3335 8188
rect 3391 8186 3415 8188
rect 3471 8186 3477 8188
rect 3231 8134 3233 8186
rect 3413 8134 3415 8186
rect 3169 8132 3175 8134
rect 3231 8132 3255 8134
rect 3311 8132 3335 8134
rect 3391 8132 3415 8134
rect 3471 8132 3477 8134
rect 3169 8123 3477 8132
rect 7608 8188 7916 8197
rect 7608 8186 7614 8188
rect 7670 8186 7694 8188
rect 7750 8186 7774 8188
rect 7830 8186 7854 8188
rect 7910 8186 7916 8188
rect 7670 8134 7672 8186
rect 7852 8134 7854 8186
rect 7608 8132 7614 8134
rect 7670 8132 7694 8134
rect 7750 8132 7774 8134
rect 7830 8132 7854 8134
rect 7910 8132 7916 8134
rect 7608 8123 7916 8132
rect 12047 8188 12355 8197
rect 12047 8186 12053 8188
rect 12109 8186 12133 8188
rect 12189 8186 12213 8188
rect 12269 8186 12293 8188
rect 12349 8186 12355 8188
rect 12109 8134 12111 8186
rect 12291 8134 12293 8186
rect 12047 8132 12053 8134
rect 12109 8132 12133 8134
rect 12189 8132 12213 8134
rect 12269 8132 12293 8134
rect 12349 8132 12355 8134
rect 12047 8123 12355 8132
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 5388 7644 5696 7653
rect 5388 7642 5394 7644
rect 5450 7642 5474 7644
rect 5530 7642 5554 7644
rect 5610 7642 5634 7644
rect 5690 7642 5696 7644
rect 5450 7590 5452 7642
rect 5632 7590 5634 7642
rect 5388 7588 5394 7590
rect 5450 7588 5474 7590
rect 5530 7588 5554 7590
rect 5610 7588 5634 7590
rect 5690 7588 5696 7590
rect 5388 7579 5696 7588
rect 9827 7644 10135 7653
rect 9827 7642 9833 7644
rect 9889 7642 9913 7644
rect 9969 7642 9993 7644
rect 10049 7642 10073 7644
rect 10129 7642 10135 7644
rect 9889 7590 9891 7642
rect 10071 7590 10073 7642
rect 9827 7588 9833 7590
rect 9889 7588 9913 7590
rect 9969 7588 9993 7590
rect 10049 7588 10073 7590
rect 10129 7588 10135 7590
rect 9827 7579 10135 7588
rect 14266 7644 14574 7653
rect 14266 7642 14272 7644
rect 14328 7642 14352 7644
rect 14408 7642 14432 7644
rect 14488 7642 14512 7644
rect 14568 7642 14574 7644
rect 14328 7590 14330 7642
rect 14510 7590 14512 7642
rect 14266 7588 14272 7590
rect 14328 7588 14352 7590
rect 14408 7588 14432 7590
rect 14488 7588 14512 7590
rect 14568 7588 14574 7590
rect 14266 7579 14574 7588
rect 14936 7546 14964 7686
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 3169 7100 3477 7109
rect 3169 7098 3175 7100
rect 3231 7098 3255 7100
rect 3311 7098 3335 7100
rect 3391 7098 3415 7100
rect 3471 7098 3477 7100
rect 3231 7046 3233 7098
rect 3413 7046 3415 7098
rect 3169 7044 3175 7046
rect 3231 7044 3255 7046
rect 3311 7044 3335 7046
rect 3391 7044 3415 7046
rect 3471 7044 3477 7046
rect 3169 7035 3477 7044
rect 7608 7100 7916 7109
rect 7608 7098 7614 7100
rect 7670 7098 7694 7100
rect 7750 7098 7774 7100
rect 7830 7098 7854 7100
rect 7910 7098 7916 7100
rect 7670 7046 7672 7098
rect 7852 7046 7854 7098
rect 7608 7044 7614 7046
rect 7670 7044 7694 7046
rect 7750 7044 7774 7046
rect 7830 7044 7854 7046
rect 7910 7044 7916 7046
rect 7608 7035 7916 7044
rect 12047 7100 12355 7109
rect 12047 7098 12053 7100
rect 12109 7098 12133 7100
rect 12189 7098 12213 7100
rect 12269 7098 12293 7100
rect 12349 7098 12355 7100
rect 12109 7046 12111 7098
rect 12291 7046 12293 7098
rect 12047 7044 12053 7046
rect 12109 7044 12133 7046
rect 12189 7044 12213 7046
rect 12269 7044 12293 7046
rect 12349 7044 12355 7046
rect 12047 7035 12355 7044
rect 15764 6866 15792 8298
rect 15948 8022 15976 8366
rect 16486 8188 16794 8197
rect 16486 8186 16492 8188
rect 16548 8186 16572 8188
rect 16628 8186 16652 8188
rect 16708 8186 16732 8188
rect 16788 8186 16794 8188
rect 16548 8134 16550 8186
rect 16730 8134 16732 8186
rect 16486 8132 16492 8134
rect 16548 8132 16572 8134
rect 16628 8132 16652 8134
rect 16708 8132 16732 8134
rect 16788 8132 16794 8134
rect 16486 8123 16794 8132
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 16396 8016 16448 8022
rect 16396 7958 16448 7964
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16132 7546 16160 7686
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 5388 6556 5696 6565
rect 5388 6554 5394 6556
rect 5450 6554 5474 6556
rect 5530 6554 5554 6556
rect 5610 6554 5634 6556
rect 5690 6554 5696 6556
rect 5450 6502 5452 6554
rect 5632 6502 5634 6554
rect 5388 6500 5394 6502
rect 5450 6500 5474 6502
rect 5530 6500 5554 6502
rect 5610 6500 5634 6502
rect 5690 6500 5696 6502
rect 5388 6491 5696 6500
rect 9827 6556 10135 6565
rect 9827 6554 9833 6556
rect 9889 6554 9913 6556
rect 9969 6554 9993 6556
rect 10049 6554 10073 6556
rect 10129 6554 10135 6556
rect 9889 6502 9891 6554
rect 10071 6502 10073 6554
rect 9827 6500 9833 6502
rect 9889 6500 9913 6502
rect 9969 6500 9993 6502
rect 10049 6500 10073 6502
rect 10129 6500 10135 6502
rect 9827 6491 10135 6500
rect 14266 6556 14574 6565
rect 14266 6554 14272 6556
rect 14328 6554 14352 6556
rect 14408 6554 14432 6556
rect 14488 6554 14512 6556
rect 14568 6554 14574 6556
rect 14328 6502 14330 6554
rect 14510 6502 14512 6554
rect 14266 6500 14272 6502
rect 14328 6500 14352 6502
rect 14408 6500 14432 6502
rect 14488 6500 14512 6502
rect 14568 6500 14574 6502
rect 14266 6491 14574 6500
rect 3169 6012 3477 6021
rect 3169 6010 3175 6012
rect 3231 6010 3255 6012
rect 3311 6010 3335 6012
rect 3391 6010 3415 6012
rect 3471 6010 3477 6012
rect 3231 5958 3233 6010
rect 3413 5958 3415 6010
rect 3169 5956 3175 5958
rect 3231 5956 3255 5958
rect 3311 5956 3335 5958
rect 3391 5956 3415 5958
rect 3471 5956 3477 5958
rect 3169 5947 3477 5956
rect 7608 6012 7916 6021
rect 7608 6010 7614 6012
rect 7670 6010 7694 6012
rect 7750 6010 7774 6012
rect 7830 6010 7854 6012
rect 7910 6010 7916 6012
rect 7670 5958 7672 6010
rect 7852 5958 7854 6010
rect 7608 5956 7614 5958
rect 7670 5956 7694 5958
rect 7750 5956 7774 5958
rect 7830 5956 7854 5958
rect 7910 5956 7916 5958
rect 7608 5947 7916 5956
rect 12047 6012 12355 6021
rect 12047 6010 12053 6012
rect 12109 6010 12133 6012
rect 12189 6010 12213 6012
rect 12269 6010 12293 6012
rect 12349 6010 12355 6012
rect 12109 5958 12111 6010
rect 12291 5958 12293 6010
rect 12047 5956 12053 5958
rect 12109 5956 12133 5958
rect 12189 5956 12213 5958
rect 12269 5956 12293 5958
rect 12349 5956 12355 5958
rect 12047 5947 12355 5956
rect 5388 5468 5696 5477
rect 5388 5466 5394 5468
rect 5450 5466 5474 5468
rect 5530 5466 5554 5468
rect 5610 5466 5634 5468
rect 5690 5466 5696 5468
rect 5450 5414 5452 5466
rect 5632 5414 5634 5466
rect 5388 5412 5394 5414
rect 5450 5412 5474 5414
rect 5530 5412 5554 5414
rect 5610 5412 5634 5414
rect 5690 5412 5696 5414
rect 5388 5403 5696 5412
rect 9827 5468 10135 5477
rect 9827 5466 9833 5468
rect 9889 5466 9913 5468
rect 9969 5466 9993 5468
rect 10049 5466 10073 5468
rect 10129 5466 10135 5468
rect 9889 5414 9891 5466
rect 10071 5414 10073 5466
rect 9827 5412 9833 5414
rect 9889 5412 9913 5414
rect 9969 5412 9993 5414
rect 10049 5412 10073 5414
rect 10129 5412 10135 5414
rect 9827 5403 10135 5412
rect 14266 5468 14574 5477
rect 14266 5466 14272 5468
rect 14328 5466 14352 5468
rect 14408 5466 14432 5468
rect 14488 5466 14512 5468
rect 14568 5466 14574 5468
rect 14328 5414 14330 5466
rect 14510 5414 14512 5466
rect 14266 5412 14272 5414
rect 14328 5412 14352 5414
rect 14408 5412 14432 5414
rect 14488 5412 14512 5414
rect 14568 5412 14574 5414
rect 14266 5403 14574 5412
rect 16040 5302 16068 6666
rect 16132 5914 16160 7142
rect 16408 7002 16436 7958
rect 16960 7954 16988 8502
rect 17052 8090 17080 28358
rect 18340 24854 18368 40326
rect 18705 40284 19013 40293
rect 18705 40282 18711 40284
rect 18767 40282 18791 40284
rect 18847 40282 18871 40284
rect 18927 40282 18951 40284
rect 19007 40282 19013 40284
rect 18767 40230 18769 40282
rect 18949 40230 18951 40282
rect 18705 40228 18711 40230
rect 18767 40228 18791 40230
rect 18847 40228 18871 40230
rect 18927 40228 18951 40230
rect 19007 40228 19013 40230
rect 18705 40219 19013 40228
rect 18705 39196 19013 39205
rect 18705 39194 18711 39196
rect 18767 39194 18791 39196
rect 18847 39194 18871 39196
rect 18927 39194 18951 39196
rect 19007 39194 19013 39196
rect 18767 39142 18769 39194
rect 18949 39142 18951 39194
rect 18705 39140 18711 39142
rect 18767 39140 18791 39142
rect 18847 39140 18871 39142
rect 18927 39140 18951 39142
rect 19007 39140 19013 39142
rect 18705 39131 19013 39140
rect 18705 38108 19013 38117
rect 18705 38106 18711 38108
rect 18767 38106 18791 38108
rect 18847 38106 18871 38108
rect 18927 38106 18951 38108
rect 19007 38106 19013 38108
rect 18767 38054 18769 38106
rect 18949 38054 18951 38106
rect 18705 38052 18711 38054
rect 18767 38052 18791 38054
rect 18847 38052 18871 38054
rect 18927 38052 18951 38054
rect 19007 38052 19013 38054
rect 18705 38043 19013 38052
rect 18705 37020 19013 37029
rect 18705 37018 18711 37020
rect 18767 37018 18791 37020
rect 18847 37018 18871 37020
rect 18927 37018 18951 37020
rect 19007 37018 19013 37020
rect 18767 36966 18769 37018
rect 18949 36966 18951 37018
rect 18705 36964 18711 36966
rect 18767 36964 18791 36966
rect 18847 36964 18871 36966
rect 18927 36964 18951 36966
rect 19007 36964 19013 36966
rect 18705 36955 19013 36964
rect 18705 35932 19013 35941
rect 18705 35930 18711 35932
rect 18767 35930 18791 35932
rect 18847 35930 18871 35932
rect 18927 35930 18951 35932
rect 19007 35930 19013 35932
rect 18767 35878 18769 35930
rect 18949 35878 18951 35930
rect 18705 35876 18711 35878
rect 18767 35876 18791 35878
rect 18847 35876 18871 35878
rect 18927 35876 18951 35878
rect 19007 35876 19013 35878
rect 18705 35867 19013 35876
rect 18705 34844 19013 34853
rect 18705 34842 18711 34844
rect 18767 34842 18791 34844
rect 18847 34842 18871 34844
rect 18927 34842 18951 34844
rect 19007 34842 19013 34844
rect 18767 34790 18769 34842
rect 18949 34790 18951 34842
rect 18705 34788 18711 34790
rect 18767 34788 18791 34790
rect 18847 34788 18871 34790
rect 18927 34788 18951 34790
rect 19007 34788 19013 34790
rect 18705 34779 19013 34788
rect 18512 34400 18564 34406
rect 18510 34368 18512 34377
rect 18564 34368 18566 34377
rect 18510 34303 18566 34312
rect 18705 33756 19013 33765
rect 18705 33754 18711 33756
rect 18767 33754 18791 33756
rect 18847 33754 18871 33756
rect 18927 33754 18951 33756
rect 19007 33754 19013 33756
rect 18767 33702 18769 33754
rect 18949 33702 18951 33754
rect 18705 33700 18711 33702
rect 18767 33700 18791 33702
rect 18847 33700 18871 33702
rect 18927 33700 18951 33702
rect 19007 33700 19013 33702
rect 18705 33691 19013 33700
rect 18705 32668 19013 32677
rect 18705 32666 18711 32668
rect 18767 32666 18791 32668
rect 18847 32666 18871 32668
rect 18927 32666 18951 32668
rect 19007 32666 19013 32668
rect 18767 32614 18769 32666
rect 18949 32614 18951 32666
rect 18705 32612 18711 32614
rect 18767 32612 18791 32614
rect 18847 32612 18871 32614
rect 18927 32612 18951 32614
rect 19007 32612 19013 32614
rect 18705 32603 19013 32612
rect 18705 31580 19013 31589
rect 18705 31578 18711 31580
rect 18767 31578 18791 31580
rect 18847 31578 18871 31580
rect 18927 31578 18951 31580
rect 19007 31578 19013 31580
rect 18767 31526 18769 31578
rect 18949 31526 18951 31578
rect 18705 31524 18711 31526
rect 18767 31524 18791 31526
rect 18847 31524 18871 31526
rect 18927 31524 18951 31526
rect 19007 31524 19013 31526
rect 18705 31515 19013 31524
rect 18705 30492 19013 30501
rect 18705 30490 18711 30492
rect 18767 30490 18791 30492
rect 18847 30490 18871 30492
rect 18927 30490 18951 30492
rect 19007 30490 19013 30492
rect 18767 30438 18769 30490
rect 18949 30438 18951 30490
rect 18705 30436 18711 30438
rect 18767 30436 18791 30438
rect 18847 30436 18871 30438
rect 18927 30436 18951 30438
rect 19007 30436 19013 30438
rect 18705 30427 19013 30436
rect 18705 29404 19013 29413
rect 18705 29402 18711 29404
rect 18767 29402 18791 29404
rect 18847 29402 18871 29404
rect 18927 29402 18951 29404
rect 19007 29402 19013 29404
rect 18767 29350 18769 29402
rect 18949 29350 18951 29402
rect 18705 29348 18711 29350
rect 18767 29348 18791 29350
rect 18847 29348 18871 29350
rect 18927 29348 18951 29350
rect 19007 29348 19013 29350
rect 18705 29339 19013 29348
rect 18604 28484 18656 28490
rect 18604 28426 18656 28432
rect 18616 28121 18644 28426
rect 18705 28316 19013 28325
rect 18705 28314 18711 28316
rect 18767 28314 18791 28316
rect 18847 28314 18871 28316
rect 18927 28314 18951 28316
rect 19007 28314 19013 28316
rect 18767 28262 18769 28314
rect 18949 28262 18951 28314
rect 18705 28260 18711 28262
rect 18767 28260 18791 28262
rect 18847 28260 18871 28262
rect 18927 28260 18951 28262
rect 19007 28260 19013 28262
rect 18705 28251 19013 28260
rect 18602 28112 18658 28121
rect 18602 28047 18658 28056
rect 18705 27228 19013 27237
rect 18705 27226 18711 27228
rect 18767 27226 18791 27228
rect 18847 27226 18871 27228
rect 18927 27226 18951 27228
rect 19007 27226 19013 27228
rect 18767 27174 18769 27226
rect 18949 27174 18951 27226
rect 18705 27172 18711 27174
rect 18767 27172 18791 27174
rect 18847 27172 18871 27174
rect 18927 27172 18951 27174
rect 19007 27172 19013 27174
rect 18705 27163 19013 27172
rect 18705 26140 19013 26149
rect 18705 26138 18711 26140
rect 18767 26138 18791 26140
rect 18847 26138 18871 26140
rect 18927 26138 18951 26140
rect 19007 26138 19013 26140
rect 18767 26086 18769 26138
rect 18949 26086 18951 26138
rect 18705 26084 18711 26086
rect 18767 26084 18791 26086
rect 18847 26084 18871 26086
rect 18927 26084 18951 26086
rect 19007 26084 19013 26086
rect 18705 26075 19013 26084
rect 18705 25052 19013 25061
rect 18705 25050 18711 25052
rect 18767 25050 18791 25052
rect 18847 25050 18871 25052
rect 18927 25050 18951 25052
rect 19007 25050 19013 25052
rect 18767 24998 18769 25050
rect 18949 24998 18951 25050
rect 18705 24996 18711 24998
rect 18767 24996 18791 24998
rect 18847 24996 18871 24998
rect 18927 24996 18951 24998
rect 19007 24996 19013 24998
rect 18705 24987 19013 24996
rect 18340 24826 18460 24854
rect 17132 16108 17184 16114
rect 17132 16050 17184 16056
rect 17144 8498 17172 16050
rect 18328 16040 18380 16046
rect 18328 15982 18380 15988
rect 18340 15609 18368 15982
rect 18326 15600 18382 15609
rect 18326 15535 18382 15544
rect 18432 8634 18460 24826
rect 18705 23964 19013 23973
rect 18705 23962 18711 23964
rect 18767 23962 18791 23964
rect 18847 23962 18871 23964
rect 18927 23962 18951 23964
rect 19007 23962 19013 23964
rect 18767 23910 18769 23962
rect 18949 23910 18951 23962
rect 18705 23908 18711 23910
rect 18767 23908 18791 23910
rect 18847 23908 18871 23910
rect 18927 23908 18951 23910
rect 19007 23908 19013 23910
rect 18705 23899 19013 23908
rect 18705 22876 19013 22885
rect 18705 22874 18711 22876
rect 18767 22874 18791 22876
rect 18847 22874 18871 22876
rect 18927 22874 18951 22876
rect 19007 22874 19013 22876
rect 18767 22822 18769 22874
rect 18949 22822 18951 22874
rect 18705 22820 18711 22822
rect 18767 22820 18791 22822
rect 18847 22820 18871 22822
rect 18927 22820 18951 22822
rect 19007 22820 19013 22822
rect 18705 22811 19013 22820
rect 18512 22228 18564 22234
rect 18512 22170 18564 22176
rect 18524 22137 18552 22170
rect 18510 22128 18566 22137
rect 18510 22063 18566 22072
rect 18705 21788 19013 21797
rect 18705 21786 18711 21788
rect 18767 21786 18791 21788
rect 18847 21786 18871 21788
rect 18927 21786 18951 21788
rect 19007 21786 19013 21788
rect 18767 21734 18769 21786
rect 18949 21734 18951 21786
rect 18705 21732 18711 21734
rect 18767 21732 18791 21734
rect 18847 21732 18871 21734
rect 18927 21732 18951 21734
rect 19007 21732 19013 21734
rect 18705 21723 19013 21732
rect 18705 20700 19013 20709
rect 18705 20698 18711 20700
rect 18767 20698 18791 20700
rect 18847 20698 18871 20700
rect 18927 20698 18951 20700
rect 19007 20698 19013 20700
rect 18767 20646 18769 20698
rect 18949 20646 18951 20698
rect 18705 20644 18711 20646
rect 18767 20644 18791 20646
rect 18847 20644 18871 20646
rect 18927 20644 18951 20646
rect 19007 20644 19013 20646
rect 18705 20635 19013 20644
rect 18705 19612 19013 19621
rect 18705 19610 18711 19612
rect 18767 19610 18791 19612
rect 18847 19610 18871 19612
rect 18927 19610 18951 19612
rect 19007 19610 19013 19612
rect 18767 19558 18769 19610
rect 18949 19558 18951 19610
rect 18705 19556 18711 19558
rect 18767 19556 18791 19558
rect 18847 19556 18871 19558
rect 18927 19556 18951 19558
rect 19007 19556 19013 19558
rect 18705 19547 19013 19556
rect 18705 18524 19013 18533
rect 18705 18522 18711 18524
rect 18767 18522 18791 18524
rect 18847 18522 18871 18524
rect 18927 18522 18951 18524
rect 19007 18522 19013 18524
rect 18767 18470 18769 18522
rect 18949 18470 18951 18522
rect 18705 18468 18711 18470
rect 18767 18468 18791 18470
rect 18847 18468 18871 18470
rect 18927 18468 18951 18470
rect 19007 18468 19013 18470
rect 18705 18459 19013 18468
rect 18705 17436 19013 17445
rect 18705 17434 18711 17436
rect 18767 17434 18791 17436
rect 18847 17434 18871 17436
rect 18927 17434 18951 17436
rect 19007 17434 19013 17436
rect 18767 17382 18769 17434
rect 18949 17382 18951 17434
rect 18705 17380 18711 17382
rect 18767 17380 18791 17382
rect 18847 17380 18871 17382
rect 18927 17380 18951 17382
rect 19007 17380 19013 17382
rect 18705 17371 19013 17380
rect 18705 16348 19013 16357
rect 18705 16346 18711 16348
rect 18767 16346 18791 16348
rect 18847 16346 18871 16348
rect 18927 16346 18951 16348
rect 19007 16346 19013 16348
rect 18767 16294 18769 16346
rect 18949 16294 18951 16346
rect 18705 16292 18711 16294
rect 18767 16292 18791 16294
rect 18847 16292 18871 16294
rect 18927 16292 18951 16294
rect 19007 16292 19013 16294
rect 18705 16283 19013 16292
rect 18705 15260 19013 15269
rect 18705 15258 18711 15260
rect 18767 15258 18791 15260
rect 18847 15258 18871 15260
rect 18927 15258 18951 15260
rect 19007 15258 19013 15260
rect 18767 15206 18769 15258
rect 18949 15206 18951 15258
rect 18705 15204 18711 15206
rect 18767 15204 18791 15206
rect 18847 15204 18871 15206
rect 18927 15204 18951 15206
rect 19007 15204 19013 15206
rect 18705 15195 19013 15204
rect 18705 14172 19013 14181
rect 18705 14170 18711 14172
rect 18767 14170 18791 14172
rect 18847 14170 18871 14172
rect 18927 14170 18951 14172
rect 19007 14170 19013 14172
rect 18767 14118 18769 14170
rect 18949 14118 18951 14170
rect 18705 14116 18711 14118
rect 18767 14116 18791 14118
rect 18847 14116 18871 14118
rect 18927 14116 18951 14118
rect 19007 14116 19013 14118
rect 18705 14107 19013 14116
rect 18705 13084 19013 13093
rect 18705 13082 18711 13084
rect 18767 13082 18791 13084
rect 18847 13082 18871 13084
rect 18927 13082 18951 13084
rect 19007 13082 19013 13084
rect 18767 13030 18769 13082
rect 18949 13030 18951 13082
rect 18705 13028 18711 13030
rect 18767 13028 18791 13030
rect 18847 13028 18871 13030
rect 18927 13028 18951 13030
rect 19007 13028 19013 13030
rect 18705 13019 19013 13028
rect 18705 11996 19013 12005
rect 18705 11994 18711 11996
rect 18767 11994 18791 11996
rect 18847 11994 18871 11996
rect 18927 11994 18951 11996
rect 19007 11994 19013 11996
rect 18767 11942 18769 11994
rect 18949 11942 18951 11994
rect 18705 11940 18711 11942
rect 18767 11940 18791 11942
rect 18847 11940 18871 11942
rect 18927 11940 18951 11942
rect 19007 11940 19013 11942
rect 18705 11931 19013 11940
rect 18705 10908 19013 10917
rect 18705 10906 18711 10908
rect 18767 10906 18791 10908
rect 18847 10906 18871 10908
rect 18927 10906 18951 10908
rect 19007 10906 19013 10908
rect 18767 10854 18769 10906
rect 18949 10854 18951 10906
rect 18705 10852 18711 10854
rect 18767 10852 18791 10854
rect 18847 10852 18871 10854
rect 18927 10852 18951 10854
rect 19007 10852 19013 10854
rect 18705 10843 19013 10852
rect 18705 9820 19013 9829
rect 18705 9818 18711 9820
rect 18767 9818 18791 9820
rect 18847 9818 18871 9820
rect 18927 9818 18951 9820
rect 19007 9818 19013 9820
rect 18767 9766 18769 9818
rect 18949 9766 18951 9818
rect 18705 9764 18711 9766
rect 18767 9764 18791 9766
rect 18847 9764 18871 9766
rect 18927 9764 18951 9766
rect 19007 9764 19013 9766
rect 18705 9755 19013 9764
rect 18512 9376 18564 9382
rect 18510 9344 18512 9353
rect 18564 9344 18566 9353
rect 18510 9279 18566 9288
rect 18705 8732 19013 8741
rect 18705 8730 18711 8732
rect 18767 8730 18791 8732
rect 18847 8730 18871 8732
rect 18927 8730 18951 8732
rect 19007 8730 19013 8732
rect 18767 8678 18769 8730
rect 18949 8678 18951 8730
rect 18705 8676 18711 8678
rect 18767 8676 18791 8678
rect 18847 8676 18871 8678
rect 18927 8676 18951 8678
rect 19007 8676 19013 8678
rect 18705 8667 19013 8676
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16776 7392 16804 7822
rect 16776 7364 16896 7392
rect 16486 7100 16794 7109
rect 16486 7098 16492 7100
rect 16548 7098 16572 7100
rect 16628 7098 16652 7100
rect 16708 7098 16732 7100
rect 16788 7098 16794 7100
rect 16548 7046 16550 7098
rect 16730 7046 16732 7098
rect 16486 7044 16492 7046
rect 16548 7044 16572 7046
rect 16628 7044 16652 7046
rect 16708 7044 16732 7046
rect 16788 7044 16794 7046
rect 16486 7035 16794 7044
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16672 6792 16724 6798
rect 16672 6734 16724 6740
rect 16684 6458 16712 6734
rect 16868 6662 16896 7364
rect 16960 6934 16988 7890
rect 16948 6928 17000 6934
rect 17144 6914 17172 8434
rect 18432 7954 18460 8570
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 17592 7744 17644 7750
rect 18144 7744 18196 7750
rect 17644 7704 17724 7732
rect 17592 7686 17644 7692
rect 17420 7002 17448 7686
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 7002 17632 7346
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 17592 6996 17644 7002
rect 17592 6938 17644 6944
rect 17696 6934 17724 7704
rect 18144 7686 18196 7692
rect 17684 6928 17736 6934
rect 17000 6886 17080 6914
rect 17144 6886 17264 6914
rect 16948 6870 17000 6876
rect 17052 6746 17080 6886
rect 17132 6792 17184 6798
rect 17052 6740 17132 6746
rect 17052 6734 17184 6740
rect 17052 6718 17172 6734
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16486 6012 16794 6021
rect 16486 6010 16492 6012
rect 16548 6010 16572 6012
rect 16628 6010 16652 6012
rect 16708 6010 16732 6012
rect 16788 6010 16794 6012
rect 16548 5958 16550 6010
rect 16730 5958 16732 6010
rect 16486 5956 16492 5958
rect 16548 5956 16572 5958
rect 16628 5956 16652 5958
rect 16708 5956 16732 5958
rect 16788 5956 16794 5958
rect 16486 5947 16794 5956
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 17052 5370 17080 6718
rect 17236 6458 17264 6886
rect 17684 6870 17736 6876
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 3169 4924 3477 4933
rect 3169 4922 3175 4924
rect 3231 4922 3255 4924
rect 3311 4922 3335 4924
rect 3391 4922 3415 4924
rect 3471 4922 3477 4924
rect 3231 4870 3233 4922
rect 3413 4870 3415 4922
rect 3169 4868 3175 4870
rect 3231 4868 3255 4870
rect 3311 4868 3335 4870
rect 3391 4868 3415 4870
rect 3471 4868 3477 4870
rect 3169 4859 3477 4868
rect 7608 4924 7916 4933
rect 7608 4922 7614 4924
rect 7670 4922 7694 4924
rect 7750 4922 7774 4924
rect 7830 4922 7854 4924
rect 7910 4922 7916 4924
rect 7670 4870 7672 4922
rect 7852 4870 7854 4922
rect 7608 4868 7614 4870
rect 7670 4868 7694 4870
rect 7750 4868 7774 4870
rect 7830 4868 7854 4870
rect 7910 4868 7916 4870
rect 7608 4859 7916 4868
rect 12047 4924 12355 4933
rect 12047 4922 12053 4924
rect 12109 4922 12133 4924
rect 12189 4922 12213 4924
rect 12269 4922 12293 4924
rect 12349 4922 12355 4924
rect 12109 4870 12111 4922
rect 12291 4870 12293 4922
rect 12047 4868 12053 4870
rect 12109 4868 12133 4870
rect 12189 4868 12213 4870
rect 12269 4868 12293 4870
rect 12349 4868 12355 4870
rect 12047 4859 12355 4868
rect 5388 4380 5696 4389
rect 5388 4378 5394 4380
rect 5450 4378 5474 4380
rect 5530 4378 5554 4380
rect 5610 4378 5634 4380
rect 5690 4378 5696 4380
rect 5450 4326 5452 4378
rect 5632 4326 5634 4378
rect 5388 4324 5394 4326
rect 5450 4324 5474 4326
rect 5530 4324 5554 4326
rect 5610 4324 5634 4326
rect 5690 4324 5696 4326
rect 5388 4315 5696 4324
rect 9827 4380 10135 4389
rect 9827 4378 9833 4380
rect 9889 4378 9913 4380
rect 9969 4378 9993 4380
rect 10049 4378 10073 4380
rect 10129 4378 10135 4380
rect 9889 4326 9891 4378
rect 10071 4326 10073 4378
rect 9827 4324 9833 4326
rect 9889 4324 9913 4326
rect 9969 4324 9993 4326
rect 10049 4324 10073 4326
rect 10129 4324 10135 4326
rect 9827 4315 10135 4324
rect 14266 4380 14574 4389
rect 14266 4378 14272 4380
rect 14328 4378 14352 4380
rect 14408 4378 14432 4380
rect 14488 4378 14512 4380
rect 14568 4378 14574 4380
rect 14328 4326 14330 4378
rect 14510 4326 14512 4378
rect 14266 4324 14272 4326
rect 14328 4324 14352 4326
rect 14408 4324 14432 4326
rect 14488 4324 14512 4326
rect 14568 4324 14574 4326
rect 14266 4315 14574 4324
rect 15948 4146 15976 4966
rect 16040 4706 16068 5238
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16040 4678 16252 4706
rect 16028 4548 16080 4554
rect 16028 4490 16080 4496
rect 16040 4282 16068 4490
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 3169 3836 3477 3845
rect 3169 3834 3175 3836
rect 3231 3834 3255 3836
rect 3311 3834 3335 3836
rect 3391 3834 3415 3836
rect 3471 3834 3477 3836
rect 3231 3782 3233 3834
rect 3413 3782 3415 3834
rect 3169 3780 3175 3782
rect 3231 3780 3255 3782
rect 3311 3780 3335 3782
rect 3391 3780 3415 3782
rect 3471 3780 3477 3782
rect 3169 3771 3477 3780
rect 7608 3836 7916 3845
rect 7608 3834 7614 3836
rect 7670 3834 7694 3836
rect 7750 3834 7774 3836
rect 7830 3834 7854 3836
rect 7910 3834 7916 3836
rect 7670 3782 7672 3834
rect 7852 3782 7854 3834
rect 7608 3780 7614 3782
rect 7670 3780 7694 3782
rect 7750 3780 7774 3782
rect 7830 3780 7854 3782
rect 7910 3780 7916 3782
rect 7608 3771 7916 3780
rect 12047 3836 12355 3845
rect 12047 3834 12053 3836
rect 12109 3834 12133 3836
rect 12189 3834 12213 3836
rect 12269 3834 12293 3836
rect 12349 3834 12355 3836
rect 12109 3782 12111 3834
rect 12291 3782 12293 3834
rect 12047 3780 12053 3782
rect 12109 3780 12133 3782
rect 12189 3780 12213 3782
rect 12269 3780 12293 3782
rect 12349 3780 12355 3782
rect 12047 3771 12355 3780
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 3169 2748 3477 2757
rect 3169 2746 3175 2748
rect 3231 2746 3255 2748
rect 3311 2746 3335 2748
rect 3391 2746 3415 2748
rect 3471 2746 3477 2748
rect 3231 2694 3233 2746
rect 3413 2694 3415 2746
rect 3169 2692 3175 2694
rect 3231 2692 3255 2694
rect 3311 2692 3335 2694
rect 3391 2692 3415 2694
rect 3471 2692 3477 2694
rect 3169 2683 3477 2692
rect 5000 800 5028 3470
rect 16132 3398 16160 4422
rect 16120 3392 16172 3398
rect 16120 3334 16172 3340
rect 5388 3292 5696 3301
rect 5388 3290 5394 3292
rect 5450 3290 5474 3292
rect 5530 3290 5554 3292
rect 5610 3290 5634 3292
rect 5690 3290 5696 3292
rect 5450 3238 5452 3290
rect 5632 3238 5634 3290
rect 5388 3236 5394 3238
rect 5450 3236 5474 3238
rect 5530 3236 5554 3238
rect 5610 3236 5634 3238
rect 5690 3236 5696 3238
rect 5388 3227 5696 3236
rect 9827 3292 10135 3301
rect 9827 3290 9833 3292
rect 9889 3290 9913 3292
rect 9969 3290 9993 3292
rect 10049 3290 10073 3292
rect 10129 3290 10135 3292
rect 9889 3238 9891 3290
rect 10071 3238 10073 3290
rect 9827 3236 9833 3238
rect 9889 3236 9913 3238
rect 9969 3236 9993 3238
rect 10049 3236 10073 3238
rect 10129 3236 10135 3238
rect 9827 3227 10135 3236
rect 14266 3292 14574 3301
rect 14266 3290 14272 3292
rect 14328 3290 14352 3292
rect 14408 3290 14432 3292
rect 14488 3290 14512 3292
rect 14568 3290 14574 3292
rect 14328 3238 14330 3290
rect 14510 3238 14512 3290
rect 14266 3236 14272 3238
rect 14328 3236 14352 3238
rect 14408 3236 14432 3238
rect 14488 3236 14512 3238
rect 14568 3236 14574 3238
rect 14266 3227 14574 3236
rect 16224 3058 16252 4678
rect 16316 4146 16344 5170
rect 16408 4146 16436 5306
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16486 4924 16794 4933
rect 16486 4922 16492 4924
rect 16548 4922 16572 4924
rect 16628 4922 16652 4924
rect 16708 4922 16732 4924
rect 16788 4922 16794 4924
rect 16548 4870 16550 4922
rect 16730 4870 16732 4922
rect 16486 4868 16492 4870
rect 16548 4868 16572 4870
rect 16628 4868 16652 4870
rect 16708 4868 16732 4870
rect 16788 4868 16794 4870
rect 16486 4859 16794 4868
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16408 3670 16436 4082
rect 16486 3836 16794 3845
rect 16486 3834 16492 3836
rect 16548 3834 16572 3836
rect 16628 3834 16652 3836
rect 16708 3834 16732 3836
rect 16788 3834 16794 3836
rect 16548 3782 16550 3834
rect 16730 3782 16732 3834
rect 16486 3780 16492 3782
rect 16548 3780 16572 3782
rect 16628 3780 16652 3782
rect 16708 3780 16732 3782
rect 16788 3780 16794 3782
rect 16486 3771 16794 3780
rect 16396 3664 16448 3670
rect 16316 3612 16396 3618
rect 16316 3606 16448 3612
rect 16316 3590 16436 3606
rect 16316 3058 16344 3590
rect 16868 3534 16896 5170
rect 17132 4480 17184 4486
rect 17236 4468 17264 6394
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5030 17448 5578
rect 17696 5166 17724 6870
rect 18156 6866 18184 7686
rect 18432 7546 18460 7890
rect 18705 7644 19013 7653
rect 18705 7642 18711 7644
rect 18767 7642 18791 7644
rect 18847 7642 18871 7644
rect 18927 7642 18951 7644
rect 19007 7642 19013 7644
rect 18767 7590 18769 7642
rect 18949 7590 18951 7642
rect 18705 7588 18711 7590
rect 18767 7588 18791 7590
rect 18847 7588 18871 7590
rect 18927 7588 18951 7590
rect 19007 7588 19013 7590
rect 18705 7579 19013 7588
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18144 6860 18196 6866
rect 18144 6802 18196 6808
rect 18705 6556 19013 6565
rect 18705 6554 18711 6556
rect 18767 6554 18791 6556
rect 18847 6554 18871 6556
rect 18927 6554 18951 6556
rect 19007 6554 19013 6556
rect 18767 6502 18769 6554
rect 18949 6502 18951 6554
rect 18705 6500 18711 6502
rect 18767 6500 18791 6502
rect 18847 6500 18871 6502
rect 18927 6500 18951 6502
rect 19007 6500 19013 6502
rect 18705 6491 19013 6500
rect 18705 5468 19013 5477
rect 18705 5466 18711 5468
rect 18767 5466 18791 5468
rect 18847 5466 18871 5468
rect 18927 5466 18951 5468
rect 19007 5466 19013 5468
rect 18767 5414 18769 5466
rect 18949 5414 18951 5466
rect 18705 5412 18711 5414
rect 18767 5412 18791 5414
rect 18847 5412 18871 5414
rect 18927 5412 18951 5414
rect 19007 5412 19013 5414
rect 18705 5403 19013 5412
rect 17684 5160 17736 5166
rect 17684 5102 17736 5108
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17316 4616 17368 4622
rect 17316 4558 17368 4564
rect 17184 4440 17264 4468
rect 17132 4422 17184 4428
rect 17144 3602 17172 4422
rect 17328 3738 17356 4558
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17420 3534 17448 4966
rect 17696 4622 17724 5102
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 18705 4380 19013 4389
rect 18705 4378 18711 4380
rect 18767 4378 18791 4380
rect 18847 4378 18871 4380
rect 18927 4378 18951 4380
rect 19007 4378 19013 4380
rect 18767 4326 18769 4378
rect 18949 4326 18951 4378
rect 18705 4324 18711 4326
rect 18767 4324 18791 4326
rect 18847 4324 18871 4326
rect 18927 4324 18951 4326
rect 19007 4324 19013 4326
rect 18705 4315 19013 4324
rect 17684 4140 17736 4146
rect 17684 4082 17736 4088
rect 16856 3528 16908 3534
rect 16856 3470 16908 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 16488 3392 16540 3398
rect 16488 3334 16540 3340
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 7608 2748 7916 2757
rect 7608 2746 7614 2748
rect 7670 2746 7694 2748
rect 7750 2746 7774 2748
rect 7830 2746 7854 2748
rect 7910 2746 7916 2748
rect 7670 2694 7672 2746
rect 7852 2694 7854 2746
rect 7608 2692 7614 2694
rect 7670 2692 7694 2694
rect 7750 2692 7774 2694
rect 7830 2692 7854 2694
rect 7910 2692 7916 2694
rect 7608 2683 7916 2692
rect 12047 2748 12355 2757
rect 12047 2746 12053 2748
rect 12109 2746 12133 2748
rect 12189 2746 12213 2748
rect 12269 2746 12293 2748
rect 12349 2746 12355 2748
rect 12109 2694 12111 2746
rect 12291 2694 12293 2746
rect 12047 2692 12053 2694
rect 12109 2692 12133 2694
rect 12189 2692 12213 2694
rect 12269 2692 12293 2694
rect 12349 2692 12355 2694
rect 12047 2683 12355 2692
rect 16224 2650 16252 2994
rect 16500 2922 16528 3334
rect 17696 3194 17724 4082
rect 18328 4072 18380 4078
rect 18328 4014 18380 4020
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 16488 2916 16540 2922
rect 16488 2858 16540 2864
rect 16486 2748 16794 2757
rect 16486 2746 16492 2748
rect 16548 2746 16572 2748
rect 16628 2746 16652 2748
rect 16708 2746 16732 2748
rect 16788 2746 16794 2748
rect 16548 2694 16550 2746
rect 16730 2694 16732 2746
rect 16486 2692 16492 2694
rect 16548 2692 16572 2694
rect 16628 2692 16652 2694
rect 16708 2692 16732 2694
rect 16788 2692 16794 2694
rect 16486 2683 16794 2692
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 17696 2514 17724 3130
rect 18340 3097 18368 4014
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18326 3088 18382 3097
rect 18326 3023 18382 3032
rect 18432 2650 18460 3402
rect 18705 3292 19013 3301
rect 18705 3290 18711 3292
rect 18767 3290 18791 3292
rect 18847 3290 18871 3292
rect 18927 3290 18951 3292
rect 19007 3290 19013 3292
rect 18767 3238 18769 3290
rect 18949 3238 18951 3290
rect 18705 3236 18711 3238
rect 18767 3236 18791 3238
rect 18847 3236 18871 3238
rect 18927 3236 18951 3238
rect 19007 3236 19013 3238
rect 18705 3227 19013 3236
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 17684 2508 17736 2514
rect 17684 2450 17736 2456
rect 15016 2440 15068 2446
rect 15016 2382 15068 2388
rect 5388 2204 5696 2213
rect 5388 2202 5394 2204
rect 5450 2202 5474 2204
rect 5530 2202 5554 2204
rect 5610 2202 5634 2204
rect 5690 2202 5696 2204
rect 5450 2150 5452 2202
rect 5632 2150 5634 2202
rect 5388 2148 5394 2150
rect 5450 2148 5474 2150
rect 5530 2148 5554 2150
rect 5610 2148 5634 2150
rect 5690 2148 5696 2150
rect 5388 2139 5696 2148
rect 9827 2204 10135 2213
rect 9827 2202 9833 2204
rect 9889 2202 9913 2204
rect 9969 2202 9993 2204
rect 10049 2202 10073 2204
rect 10129 2202 10135 2204
rect 9889 2150 9891 2202
rect 10071 2150 10073 2202
rect 9827 2148 9833 2150
rect 9889 2148 9913 2150
rect 9969 2148 9993 2150
rect 10049 2148 10073 2150
rect 10129 2148 10135 2150
rect 9827 2139 10135 2148
rect 14266 2204 14574 2213
rect 14266 2202 14272 2204
rect 14328 2202 14352 2204
rect 14408 2202 14432 2204
rect 14488 2202 14512 2204
rect 14568 2202 14574 2204
rect 14328 2150 14330 2202
rect 14510 2150 14512 2202
rect 14266 2148 14272 2150
rect 14328 2148 14352 2150
rect 14408 2148 14432 2150
rect 14488 2148 14512 2150
rect 14568 2148 14574 2150
rect 14266 2139 14574 2148
rect 15028 1306 15056 2382
rect 18705 2204 19013 2213
rect 18705 2202 18711 2204
rect 18767 2202 18791 2204
rect 18847 2202 18871 2204
rect 18927 2202 18951 2204
rect 19007 2202 19013 2204
rect 18767 2150 18769 2202
rect 18949 2150 18951 2202
rect 18705 2148 18711 2150
rect 18767 2148 18791 2150
rect 18847 2148 18871 2150
rect 18927 2148 18951 2150
rect 19007 2148 19013 2150
rect 18705 2139 19013 2148
rect 14936 1278 15056 1306
rect 14936 800 14964 1278
rect 4986 0 5042 800
rect 14922 0 14978 800
<< via2 >>
rect 3175 47354 3231 47356
rect 3255 47354 3311 47356
rect 3335 47354 3391 47356
rect 3415 47354 3471 47356
rect 3175 47302 3221 47354
rect 3221 47302 3231 47354
rect 3255 47302 3285 47354
rect 3285 47302 3297 47354
rect 3297 47302 3311 47354
rect 3335 47302 3349 47354
rect 3349 47302 3361 47354
rect 3361 47302 3391 47354
rect 3415 47302 3425 47354
rect 3425 47302 3471 47354
rect 3175 47300 3231 47302
rect 3255 47300 3311 47302
rect 3335 47300 3391 47302
rect 3415 47300 3471 47302
rect 7614 47354 7670 47356
rect 7694 47354 7750 47356
rect 7774 47354 7830 47356
rect 7854 47354 7910 47356
rect 7614 47302 7660 47354
rect 7660 47302 7670 47354
rect 7694 47302 7724 47354
rect 7724 47302 7736 47354
rect 7736 47302 7750 47354
rect 7774 47302 7788 47354
rect 7788 47302 7800 47354
rect 7800 47302 7830 47354
rect 7854 47302 7864 47354
rect 7864 47302 7910 47354
rect 7614 47300 7670 47302
rect 7694 47300 7750 47302
rect 7774 47300 7830 47302
rect 7854 47300 7910 47302
rect 12053 47354 12109 47356
rect 12133 47354 12189 47356
rect 12213 47354 12269 47356
rect 12293 47354 12349 47356
rect 12053 47302 12099 47354
rect 12099 47302 12109 47354
rect 12133 47302 12163 47354
rect 12163 47302 12175 47354
rect 12175 47302 12189 47354
rect 12213 47302 12227 47354
rect 12227 47302 12239 47354
rect 12239 47302 12269 47354
rect 12293 47302 12303 47354
rect 12303 47302 12349 47354
rect 12053 47300 12109 47302
rect 12133 47300 12189 47302
rect 12213 47300 12269 47302
rect 12293 47300 12349 47302
rect 16492 47354 16548 47356
rect 16572 47354 16628 47356
rect 16652 47354 16708 47356
rect 16732 47354 16788 47356
rect 16492 47302 16538 47354
rect 16538 47302 16548 47354
rect 16572 47302 16602 47354
rect 16602 47302 16614 47354
rect 16614 47302 16628 47354
rect 16652 47302 16666 47354
rect 16666 47302 16678 47354
rect 16678 47302 16708 47354
rect 16732 47302 16742 47354
rect 16742 47302 16788 47354
rect 16492 47300 16548 47302
rect 16572 47300 16628 47302
rect 16652 47300 16708 47302
rect 16732 47300 16788 47302
rect 18510 47096 18566 47152
rect 5394 46810 5450 46812
rect 5474 46810 5530 46812
rect 5554 46810 5610 46812
rect 5634 46810 5690 46812
rect 5394 46758 5440 46810
rect 5440 46758 5450 46810
rect 5474 46758 5504 46810
rect 5504 46758 5516 46810
rect 5516 46758 5530 46810
rect 5554 46758 5568 46810
rect 5568 46758 5580 46810
rect 5580 46758 5610 46810
rect 5634 46758 5644 46810
rect 5644 46758 5690 46810
rect 5394 46756 5450 46758
rect 5474 46756 5530 46758
rect 5554 46756 5610 46758
rect 5634 46756 5690 46758
rect 9833 46810 9889 46812
rect 9913 46810 9969 46812
rect 9993 46810 10049 46812
rect 10073 46810 10129 46812
rect 9833 46758 9879 46810
rect 9879 46758 9889 46810
rect 9913 46758 9943 46810
rect 9943 46758 9955 46810
rect 9955 46758 9969 46810
rect 9993 46758 10007 46810
rect 10007 46758 10019 46810
rect 10019 46758 10049 46810
rect 10073 46758 10083 46810
rect 10083 46758 10129 46810
rect 9833 46756 9889 46758
rect 9913 46756 9969 46758
rect 9993 46756 10049 46758
rect 10073 46756 10129 46758
rect 14272 46810 14328 46812
rect 14352 46810 14408 46812
rect 14432 46810 14488 46812
rect 14512 46810 14568 46812
rect 14272 46758 14318 46810
rect 14318 46758 14328 46810
rect 14352 46758 14382 46810
rect 14382 46758 14394 46810
rect 14394 46758 14408 46810
rect 14432 46758 14446 46810
rect 14446 46758 14458 46810
rect 14458 46758 14488 46810
rect 14512 46758 14522 46810
rect 14522 46758 14568 46810
rect 14272 46756 14328 46758
rect 14352 46756 14408 46758
rect 14432 46756 14488 46758
rect 14512 46756 14568 46758
rect 18711 46810 18767 46812
rect 18791 46810 18847 46812
rect 18871 46810 18927 46812
rect 18951 46810 19007 46812
rect 18711 46758 18757 46810
rect 18757 46758 18767 46810
rect 18791 46758 18821 46810
rect 18821 46758 18833 46810
rect 18833 46758 18847 46810
rect 18871 46758 18885 46810
rect 18885 46758 18897 46810
rect 18897 46758 18927 46810
rect 18951 46758 18961 46810
rect 18961 46758 19007 46810
rect 18711 46756 18767 46758
rect 18791 46756 18847 46758
rect 18871 46756 18927 46758
rect 18951 46756 19007 46758
rect 3175 46266 3231 46268
rect 3255 46266 3311 46268
rect 3335 46266 3391 46268
rect 3415 46266 3471 46268
rect 3175 46214 3221 46266
rect 3221 46214 3231 46266
rect 3255 46214 3285 46266
rect 3285 46214 3297 46266
rect 3297 46214 3311 46266
rect 3335 46214 3349 46266
rect 3349 46214 3361 46266
rect 3361 46214 3391 46266
rect 3415 46214 3425 46266
rect 3425 46214 3471 46266
rect 3175 46212 3231 46214
rect 3255 46212 3311 46214
rect 3335 46212 3391 46214
rect 3415 46212 3471 46214
rect 7614 46266 7670 46268
rect 7694 46266 7750 46268
rect 7774 46266 7830 46268
rect 7854 46266 7910 46268
rect 7614 46214 7660 46266
rect 7660 46214 7670 46266
rect 7694 46214 7724 46266
rect 7724 46214 7736 46266
rect 7736 46214 7750 46266
rect 7774 46214 7788 46266
rect 7788 46214 7800 46266
rect 7800 46214 7830 46266
rect 7854 46214 7864 46266
rect 7864 46214 7910 46266
rect 7614 46212 7670 46214
rect 7694 46212 7750 46214
rect 7774 46212 7830 46214
rect 7854 46212 7910 46214
rect 12053 46266 12109 46268
rect 12133 46266 12189 46268
rect 12213 46266 12269 46268
rect 12293 46266 12349 46268
rect 12053 46214 12099 46266
rect 12099 46214 12109 46266
rect 12133 46214 12163 46266
rect 12163 46214 12175 46266
rect 12175 46214 12189 46266
rect 12213 46214 12227 46266
rect 12227 46214 12239 46266
rect 12239 46214 12269 46266
rect 12293 46214 12303 46266
rect 12303 46214 12349 46266
rect 12053 46212 12109 46214
rect 12133 46212 12189 46214
rect 12213 46212 12269 46214
rect 12293 46212 12349 46214
rect 16492 46266 16548 46268
rect 16572 46266 16628 46268
rect 16652 46266 16708 46268
rect 16732 46266 16788 46268
rect 16492 46214 16538 46266
rect 16538 46214 16548 46266
rect 16572 46214 16602 46266
rect 16602 46214 16614 46266
rect 16614 46214 16628 46266
rect 16652 46214 16666 46266
rect 16666 46214 16678 46266
rect 16678 46214 16708 46266
rect 16732 46214 16742 46266
rect 16742 46214 16788 46266
rect 16492 46212 16548 46214
rect 16572 46212 16628 46214
rect 16652 46212 16708 46214
rect 16732 46212 16788 46214
rect 5394 45722 5450 45724
rect 5474 45722 5530 45724
rect 5554 45722 5610 45724
rect 5634 45722 5690 45724
rect 5394 45670 5440 45722
rect 5440 45670 5450 45722
rect 5474 45670 5504 45722
rect 5504 45670 5516 45722
rect 5516 45670 5530 45722
rect 5554 45670 5568 45722
rect 5568 45670 5580 45722
rect 5580 45670 5610 45722
rect 5634 45670 5644 45722
rect 5644 45670 5690 45722
rect 5394 45668 5450 45670
rect 5474 45668 5530 45670
rect 5554 45668 5610 45670
rect 5634 45668 5690 45670
rect 9833 45722 9889 45724
rect 9913 45722 9969 45724
rect 9993 45722 10049 45724
rect 10073 45722 10129 45724
rect 9833 45670 9879 45722
rect 9879 45670 9889 45722
rect 9913 45670 9943 45722
rect 9943 45670 9955 45722
rect 9955 45670 9969 45722
rect 9993 45670 10007 45722
rect 10007 45670 10019 45722
rect 10019 45670 10049 45722
rect 10073 45670 10083 45722
rect 10083 45670 10129 45722
rect 9833 45668 9889 45670
rect 9913 45668 9969 45670
rect 9993 45668 10049 45670
rect 10073 45668 10129 45670
rect 14272 45722 14328 45724
rect 14352 45722 14408 45724
rect 14432 45722 14488 45724
rect 14512 45722 14568 45724
rect 14272 45670 14318 45722
rect 14318 45670 14328 45722
rect 14352 45670 14382 45722
rect 14382 45670 14394 45722
rect 14394 45670 14408 45722
rect 14432 45670 14446 45722
rect 14446 45670 14458 45722
rect 14458 45670 14488 45722
rect 14512 45670 14522 45722
rect 14522 45670 14568 45722
rect 14272 45668 14328 45670
rect 14352 45668 14408 45670
rect 14432 45668 14488 45670
rect 14512 45668 14568 45670
rect 18711 45722 18767 45724
rect 18791 45722 18847 45724
rect 18871 45722 18927 45724
rect 18951 45722 19007 45724
rect 18711 45670 18757 45722
rect 18757 45670 18767 45722
rect 18791 45670 18821 45722
rect 18821 45670 18833 45722
rect 18833 45670 18847 45722
rect 18871 45670 18885 45722
rect 18885 45670 18897 45722
rect 18897 45670 18927 45722
rect 18951 45670 18961 45722
rect 18961 45670 19007 45722
rect 18711 45668 18767 45670
rect 18791 45668 18847 45670
rect 18871 45668 18927 45670
rect 18951 45668 19007 45670
rect 3175 45178 3231 45180
rect 3255 45178 3311 45180
rect 3335 45178 3391 45180
rect 3415 45178 3471 45180
rect 3175 45126 3221 45178
rect 3221 45126 3231 45178
rect 3255 45126 3285 45178
rect 3285 45126 3297 45178
rect 3297 45126 3311 45178
rect 3335 45126 3349 45178
rect 3349 45126 3361 45178
rect 3361 45126 3391 45178
rect 3415 45126 3425 45178
rect 3425 45126 3471 45178
rect 3175 45124 3231 45126
rect 3255 45124 3311 45126
rect 3335 45124 3391 45126
rect 3415 45124 3471 45126
rect 7614 45178 7670 45180
rect 7694 45178 7750 45180
rect 7774 45178 7830 45180
rect 7854 45178 7910 45180
rect 7614 45126 7660 45178
rect 7660 45126 7670 45178
rect 7694 45126 7724 45178
rect 7724 45126 7736 45178
rect 7736 45126 7750 45178
rect 7774 45126 7788 45178
rect 7788 45126 7800 45178
rect 7800 45126 7830 45178
rect 7854 45126 7864 45178
rect 7864 45126 7910 45178
rect 7614 45124 7670 45126
rect 7694 45124 7750 45126
rect 7774 45124 7830 45126
rect 7854 45124 7910 45126
rect 12053 45178 12109 45180
rect 12133 45178 12189 45180
rect 12213 45178 12269 45180
rect 12293 45178 12349 45180
rect 12053 45126 12099 45178
rect 12099 45126 12109 45178
rect 12133 45126 12163 45178
rect 12163 45126 12175 45178
rect 12175 45126 12189 45178
rect 12213 45126 12227 45178
rect 12227 45126 12239 45178
rect 12239 45126 12269 45178
rect 12293 45126 12303 45178
rect 12303 45126 12349 45178
rect 12053 45124 12109 45126
rect 12133 45124 12189 45126
rect 12213 45124 12269 45126
rect 12293 45124 12349 45126
rect 16492 45178 16548 45180
rect 16572 45178 16628 45180
rect 16652 45178 16708 45180
rect 16732 45178 16788 45180
rect 16492 45126 16538 45178
rect 16538 45126 16548 45178
rect 16572 45126 16602 45178
rect 16602 45126 16614 45178
rect 16614 45126 16628 45178
rect 16652 45126 16666 45178
rect 16666 45126 16678 45178
rect 16678 45126 16708 45178
rect 16732 45126 16742 45178
rect 16742 45126 16788 45178
rect 16492 45124 16548 45126
rect 16572 45124 16628 45126
rect 16652 45124 16708 45126
rect 16732 45124 16788 45126
rect 5394 44634 5450 44636
rect 5474 44634 5530 44636
rect 5554 44634 5610 44636
rect 5634 44634 5690 44636
rect 5394 44582 5440 44634
rect 5440 44582 5450 44634
rect 5474 44582 5504 44634
rect 5504 44582 5516 44634
rect 5516 44582 5530 44634
rect 5554 44582 5568 44634
rect 5568 44582 5580 44634
rect 5580 44582 5610 44634
rect 5634 44582 5644 44634
rect 5644 44582 5690 44634
rect 5394 44580 5450 44582
rect 5474 44580 5530 44582
rect 5554 44580 5610 44582
rect 5634 44580 5690 44582
rect 9833 44634 9889 44636
rect 9913 44634 9969 44636
rect 9993 44634 10049 44636
rect 10073 44634 10129 44636
rect 9833 44582 9879 44634
rect 9879 44582 9889 44634
rect 9913 44582 9943 44634
rect 9943 44582 9955 44634
rect 9955 44582 9969 44634
rect 9993 44582 10007 44634
rect 10007 44582 10019 44634
rect 10019 44582 10049 44634
rect 10073 44582 10083 44634
rect 10083 44582 10129 44634
rect 9833 44580 9889 44582
rect 9913 44580 9969 44582
rect 9993 44580 10049 44582
rect 10073 44580 10129 44582
rect 14272 44634 14328 44636
rect 14352 44634 14408 44636
rect 14432 44634 14488 44636
rect 14512 44634 14568 44636
rect 14272 44582 14318 44634
rect 14318 44582 14328 44634
rect 14352 44582 14382 44634
rect 14382 44582 14394 44634
rect 14394 44582 14408 44634
rect 14432 44582 14446 44634
rect 14446 44582 14458 44634
rect 14458 44582 14488 44634
rect 14512 44582 14522 44634
rect 14522 44582 14568 44634
rect 14272 44580 14328 44582
rect 14352 44580 14408 44582
rect 14432 44580 14488 44582
rect 14512 44580 14568 44582
rect 18711 44634 18767 44636
rect 18791 44634 18847 44636
rect 18871 44634 18927 44636
rect 18951 44634 19007 44636
rect 18711 44582 18757 44634
rect 18757 44582 18767 44634
rect 18791 44582 18821 44634
rect 18821 44582 18833 44634
rect 18833 44582 18847 44634
rect 18871 44582 18885 44634
rect 18885 44582 18897 44634
rect 18897 44582 18927 44634
rect 18951 44582 18961 44634
rect 18961 44582 19007 44634
rect 18711 44580 18767 44582
rect 18791 44580 18847 44582
rect 18871 44580 18927 44582
rect 18951 44580 19007 44582
rect 3175 44090 3231 44092
rect 3255 44090 3311 44092
rect 3335 44090 3391 44092
rect 3415 44090 3471 44092
rect 3175 44038 3221 44090
rect 3221 44038 3231 44090
rect 3255 44038 3285 44090
rect 3285 44038 3297 44090
rect 3297 44038 3311 44090
rect 3335 44038 3349 44090
rect 3349 44038 3361 44090
rect 3361 44038 3391 44090
rect 3415 44038 3425 44090
rect 3425 44038 3471 44090
rect 3175 44036 3231 44038
rect 3255 44036 3311 44038
rect 3335 44036 3391 44038
rect 3415 44036 3471 44038
rect 7614 44090 7670 44092
rect 7694 44090 7750 44092
rect 7774 44090 7830 44092
rect 7854 44090 7910 44092
rect 7614 44038 7660 44090
rect 7660 44038 7670 44090
rect 7694 44038 7724 44090
rect 7724 44038 7736 44090
rect 7736 44038 7750 44090
rect 7774 44038 7788 44090
rect 7788 44038 7800 44090
rect 7800 44038 7830 44090
rect 7854 44038 7864 44090
rect 7864 44038 7910 44090
rect 7614 44036 7670 44038
rect 7694 44036 7750 44038
rect 7774 44036 7830 44038
rect 7854 44036 7910 44038
rect 12053 44090 12109 44092
rect 12133 44090 12189 44092
rect 12213 44090 12269 44092
rect 12293 44090 12349 44092
rect 12053 44038 12099 44090
rect 12099 44038 12109 44090
rect 12133 44038 12163 44090
rect 12163 44038 12175 44090
rect 12175 44038 12189 44090
rect 12213 44038 12227 44090
rect 12227 44038 12239 44090
rect 12239 44038 12269 44090
rect 12293 44038 12303 44090
rect 12303 44038 12349 44090
rect 12053 44036 12109 44038
rect 12133 44036 12189 44038
rect 12213 44036 12269 44038
rect 12293 44036 12349 44038
rect 16492 44090 16548 44092
rect 16572 44090 16628 44092
rect 16652 44090 16708 44092
rect 16732 44090 16788 44092
rect 16492 44038 16538 44090
rect 16538 44038 16548 44090
rect 16572 44038 16602 44090
rect 16602 44038 16614 44090
rect 16614 44038 16628 44090
rect 16652 44038 16666 44090
rect 16666 44038 16678 44090
rect 16678 44038 16708 44090
rect 16732 44038 16742 44090
rect 16742 44038 16788 44090
rect 16492 44036 16548 44038
rect 16572 44036 16628 44038
rect 16652 44036 16708 44038
rect 16732 44036 16788 44038
rect 5394 43546 5450 43548
rect 5474 43546 5530 43548
rect 5554 43546 5610 43548
rect 5634 43546 5690 43548
rect 5394 43494 5440 43546
rect 5440 43494 5450 43546
rect 5474 43494 5504 43546
rect 5504 43494 5516 43546
rect 5516 43494 5530 43546
rect 5554 43494 5568 43546
rect 5568 43494 5580 43546
rect 5580 43494 5610 43546
rect 5634 43494 5644 43546
rect 5644 43494 5690 43546
rect 5394 43492 5450 43494
rect 5474 43492 5530 43494
rect 5554 43492 5610 43494
rect 5634 43492 5690 43494
rect 9833 43546 9889 43548
rect 9913 43546 9969 43548
rect 9993 43546 10049 43548
rect 10073 43546 10129 43548
rect 9833 43494 9879 43546
rect 9879 43494 9889 43546
rect 9913 43494 9943 43546
rect 9943 43494 9955 43546
rect 9955 43494 9969 43546
rect 9993 43494 10007 43546
rect 10007 43494 10019 43546
rect 10019 43494 10049 43546
rect 10073 43494 10083 43546
rect 10083 43494 10129 43546
rect 9833 43492 9889 43494
rect 9913 43492 9969 43494
rect 9993 43492 10049 43494
rect 10073 43492 10129 43494
rect 14272 43546 14328 43548
rect 14352 43546 14408 43548
rect 14432 43546 14488 43548
rect 14512 43546 14568 43548
rect 14272 43494 14318 43546
rect 14318 43494 14328 43546
rect 14352 43494 14382 43546
rect 14382 43494 14394 43546
rect 14394 43494 14408 43546
rect 14432 43494 14446 43546
rect 14446 43494 14458 43546
rect 14458 43494 14488 43546
rect 14512 43494 14522 43546
rect 14522 43494 14568 43546
rect 14272 43492 14328 43494
rect 14352 43492 14408 43494
rect 14432 43492 14488 43494
rect 14512 43492 14568 43494
rect 18711 43546 18767 43548
rect 18791 43546 18847 43548
rect 18871 43546 18927 43548
rect 18951 43546 19007 43548
rect 18711 43494 18757 43546
rect 18757 43494 18767 43546
rect 18791 43494 18821 43546
rect 18821 43494 18833 43546
rect 18833 43494 18847 43546
rect 18871 43494 18885 43546
rect 18885 43494 18897 43546
rect 18897 43494 18927 43546
rect 18951 43494 18961 43546
rect 18961 43494 19007 43546
rect 18711 43492 18767 43494
rect 18791 43492 18847 43494
rect 18871 43492 18927 43494
rect 18951 43492 19007 43494
rect 3175 43002 3231 43004
rect 3255 43002 3311 43004
rect 3335 43002 3391 43004
rect 3415 43002 3471 43004
rect 3175 42950 3221 43002
rect 3221 42950 3231 43002
rect 3255 42950 3285 43002
rect 3285 42950 3297 43002
rect 3297 42950 3311 43002
rect 3335 42950 3349 43002
rect 3349 42950 3361 43002
rect 3361 42950 3391 43002
rect 3415 42950 3425 43002
rect 3425 42950 3471 43002
rect 3175 42948 3231 42950
rect 3255 42948 3311 42950
rect 3335 42948 3391 42950
rect 3415 42948 3471 42950
rect 7614 43002 7670 43004
rect 7694 43002 7750 43004
rect 7774 43002 7830 43004
rect 7854 43002 7910 43004
rect 7614 42950 7660 43002
rect 7660 42950 7670 43002
rect 7694 42950 7724 43002
rect 7724 42950 7736 43002
rect 7736 42950 7750 43002
rect 7774 42950 7788 43002
rect 7788 42950 7800 43002
rect 7800 42950 7830 43002
rect 7854 42950 7864 43002
rect 7864 42950 7910 43002
rect 7614 42948 7670 42950
rect 7694 42948 7750 42950
rect 7774 42948 7830 42950
rect 7854 42948 7910 42950
rect 12053 43002 12109 43004
rect 12133 43002 12189 43004
rect 12213 43002 12269 43004
rect 12293 43002 12349 43004
rect 12053 42950 12099 43002
rect 12099 42950 12109 43002
rect 12133 42950 12163 43002
rect 12163 42950 12175 43002
rect 12175 42950 12189 43002
rect 12213 42950 12227 43002
rect 12227 42950 12239 43002
rect 12239 42950 12269 43002
rect 12293 42950 12303 43002
rect 12303 42950 12349 43002
rect 12053 42948 12109 42950
rect 12133 42948 12189 42950
rect 12213 42948 12269 42950
rect 12293 42948 12349 42950
rect 16492 43002 16548 43004
rect 16572 43002 16628 43004
rect 16652 43002 16708 43004
rect 16732 43002 16788 43004
rect 16492 42950 16538 43002
rect 16538 42950 16548 43002
rect 16572 42950 16602 43002
rect 16602 42950 16614 43002
rect 16614 42950 16628 43002
rect 16652 42950 16666 43002
rect 16666 42950 16678 43002
rect 16678 42950 16708 43002
rect 16732 42950 16742 43002
rect 16742 42950 16788 43002
rect 16492 42948 16548 42950
rect 16572 42948 16628 42950
rect 16652 42948 16708 42950
rect 16732 42948 16788 42950
rect 5394 42458 5450 42460
rect 5474 42458 5530 42460
rect 5554 42458 5610 42460
rect 5634 42458 5690 42460
rect 5394 42406 5440 42458
rect 5440 42406 5450 42458
rect 5474 42406 5504 42458
rect 5504 42406 5516 42458
rect 5516 42406 5530 42458
rect 5554 42406 5568 42458
rect 5568 42406 5580 42458
rect 5580 42406 5610 42458
rect 5634 42406 5644 42458
rect 5644 42406 5690 42458
rect 5394 42404 5450 42406
rect 5474 42404 5530 42406
rect 5554 42404 5610 42406
rect 5634 42404 5690 42406
rect 9833 42458 9889 42460
rect 9913 42458 9969 42460
rect 9993 42458 10049 42460
rect 10073 42458 10129 42460
rect 9833 42406 9879 42458
rect 9879 42406 9889 42458
rect 9913 42406 9943 42458
rect 9943 42406 9955 42458
rect 9955 42406 9969 42458
rect 9993 42406 10007 42458
rect 10007 42406 10019 42458
rect 10019 42406 10049 42458
rect 10073 42406 10083 42458
rect 10083 42406 10129 42458
rect 9833 42404 9889 42406
rect 9913 42404 9969 42406
rect 9993 42404 10049 42406
rect 10073 42404 10129 42406
rect 14272 42458 14328 42460
rect 14352 42458 14408 42460
rect 14432 42458 14488 42460
rect 14512 42458 14568 42460
rect 14272 42406 14318 42458
rect 14318 42406 14328 42458
rect 14352 42406 14382 42458
rect 14382 42406 14394 42458
rect 14394 42406 14408 42458
rect 14432 42406 14446 42458
rect 14446 42406 14458 42458
rect 14458 42406 14488 42458
rect 14512 42406 14522 42458
rect 14522 42406 14568 42458
rect 14272 42404 14328 42406
rect 14352 42404 14408 42406
rect 14432 42404 14488 42406
rect 14512 42404 14568 42406
rect 18711 42458 18767 42460
rect 18791 42458 18847 42460
rect 18871 42458 18927 42460
rect 18951 42458 19007 42460
rect 18711 42406 18757 42458
rect 18757 42406 18767 42458
rect 18791 42406 18821 42458
rect 18821 42406 18833 42458
rect 18833 42406 18847 42458
rect 18871 42406 18885 42458
rect 18885 42406 18897 42458
rect 18897 42406 18927 42458
rect 18951 42406 18961 42458
rect 18961 42406 19007 42458
rect 18711 42404 18767 42406
rect 18791 42404 18847 42406
rect 18871 42404 18927 42406
rect 18951 42404 19007 42406
rect 3175 41914 3231 41916
rect 3255 41914 3311 41916
rect 3335 41914 3391 41916
rect 3415 41914 3471 41916
rect 3175 41862 3221 41914
rect 3221 41862 3231 41914
rect 3255 41862 3285 41914
rect 3285 41862 3297 41914
rect 3297 41862 3311 41914
rect 3335 41862 3349 41914
rect 3349 41862 3361 41914
rect 3361 41862 3391 41914
rect 3415 41862 3425 41914
rect 3425 41862 3471 41914
rect 3175 41860 3231 41862
rect 3255 41860 3311 41862
rect 3335 41860 3391 41862
rect 3415 41860 3471 41862
rect 7614 41914 7670 41916
rect 7694 41914 7750 41916
rect 7774 41914 7830 41916
rect 7854 41914 7910 41916
rect 7614 41862 7660 41914
rect 7660 41862 7670 41914
rect 7694 41862 7724 41914
rect 7724 41862 7736 41914
rect 7736 41862 7750 41914
rect 7774 41862 7788 41914
rect 7788 41862 7800 41914
rect 7800 41862 7830 41914
rect 7854 41862 7864 41914
rect 7864 41862 7910 41914
rect 7614 41860 7670 41862
rect 7694 41860 7750 41862
rect 7774 41860 7830 41862
rect 7854 41860 7910 41862
rect 12053 41914 12109 41916
rect 12133 41914 12189 41916
rect 12213 41914 12269 41916
rect 12293 41914 12349 41916
rect 12053 41862 12099 41914
rect 12099 41862 12109 41914
rect 12133 41862 12163 41914
rect 12163 41862 12175 41914
rect 12175 41862 12189 41914
rect 12213 41862 12227 41914
rect 12227 41862 12239 41914
rect 12239 41862 12269 41914
rect 12293 41862 12303 41914
rect 12303 41862 12349 41914
rect 12053 41860 12109 41862
rect 12133 41860 12189 41862
rect 12213 41860 12269 41862
rect 12293 41860 12349 41862
rect 16492 41914 16548 41916
rect 16572 41914 16628 41916
rect 16652 41914 16708 41916
rect 16732 41914 16788 41916
rect 16492 41862 16538 41914
rect 16538 41862 16548 41914
rect 16572 41862 16602 41914
rect 16602 41862 16614 41914
rect 16614 41862 16628 41914
rect 16652 41862 16666 41914
rect 16666 41862 16678 41914
rect 16678 41862 16708 41914
rect 16732 41862 16742 41914
rect 16742 41862 16788 41914
rect 16492 41860 16548 41862
rect 16572 41860 16628 41862
rect 16652 41860 16708 41862
rect 16732 41860 16788 41862
rect 5394 41370 5450 41372
rect 5474 41370 5530 41372
rect 5554 41370 5610 41372
rect 5634 41370 5690 41372
rect 5394 41318 5440 41370
rect 5440 41318 5450 41370
rect 5474 41318 5504 41370
rect 5504 41318 5516 41370
rect 5516 41318 5530 41370
rect 5554 41318 5568 41370
rect 5568 41318 5580 41370
rect 5580 41318 5610 41370
rect 5634 41318 5644 41370
rect 5644 41318 5690 41370
rect 5394 41316 5450 41318
rect 5474 41316 5530 41318
rect 5554 41316 5610 41318
rect 5634 41316 5690 41318
rect 9833 41370 9889 41372
rect 9913 41370 9969 41372
rect 9993 41370 10049 41372
rect 10073 41370 10129 41372
rect 9833 41318 9879 41370
rect 9879 41318 9889 41370
rect 9913 41318 9943 41370
rect 9943 41318 9955 41370
rect 9955 41318 9969 41370
rect 9993 41318 10007 41370
rect 10007 41318 10019 41370
rect 10019 41318 10049 41370
rect 10073 41318 10083 41370
rect 10083 41318 10129 41370
rect 9833 41316 9889 41318
rect 9913 41316 9969 41318
rect 9993 41316 10049 41318
rect 10073 41316 10129 41318
rect 14272 41370 14328 41372
rect 14352 41370 14408 41372
rect 14432 41370 14488 41372
rect 14512 41370 14568 41372
rect 14272 41318 14318 41370
rect 14318 41318 14328 41370
rect 14352 41318 14382 41370
rect 14382 41318 14394 41370
rect 14394 41318 14408 41370
rect 14432 41318 14446 41370
rect 14446 41318 14458 41370
rect 14458 41318 14488 41370
rect 14512 41318 14522 41370
rect 14522 41318 14568 41370
rect 14272 41316 14328 41318
rect 14352 41316 14408 41318
rect 14432 41316 14488 41318
rect 14512 41316 14568 41318
rect 18711 41370 18767 41372
rect 18791 41370 18847 41372
rect 18871 41370 18927 41372
rect 18951 41370 19007 41372
rect 18711 41318 18757 41370
rect 18757 41318 18767 41370
rect 18791 41318 18821 41370
rect 18821 41318 18833 41370
rect 18833 41318 18847 41370
rect 18871 41318 18885 41370
rect 18885 41318 18897 41370
rect 18897 41318 18927 41370
rect 18951 41318 18961 41370
rect 18961 41318 19007 41370
rect 18711 41316 18767 41318
rect 18791 41316 18847 41318
rect 18871 41316 18927 41318
rect 18951 41316 19007 41318
rect 3175 40826 3231 40828
rect 3255 40826 3311 40828
rect 3335 40826 3391 40828
rect 3415 40826 3471 40828
rect 3175 40774 3221 40826
rect 3221 40774 3231 40826
rect 3255 40774 3285 40826
rect 3285 40774 3297 40826
rect 3297 40774 3311 40826
rect 3335 40774 3349 40826
rect 3349 40774 3361 40826
rect 3361 40774 3391 40826
rect 3415 40774 3425 40826
rect 3425 40774 3471 40826
rect 3175 40772 3231 40774
rect 3255 40772 3311 40774
rect 3335 40772 3391 40774
rect 3415 40772 3471 40774
rect 7614 40826 7670 40828
rect 7694 40826 7750 40828
rect 7774 40826 7830 40828
rect 7854 40826 7910 40828
rect 7614 40774 7660 40826
rect 7660 40774 7670 40826
rect 7694 40774 7724 40826
rect 7724 40774 7736 40826
rect 7736 40774 7750 40826
rect 7774 40774 7788 40826
rect 7788 40774 7800 40826
rect 7800 40774 7830 40826
rect 7854 40774 7864 40826
rect 7864 40774 7910 40826
rect 7614 40772 7670 40774
rect 7694 40772 7750 40774
rect 7774 40772 7830 40774
rect 7854 40772 7910 40774
rect 12053 40826 12109 40828
rect 12133 40826 12189 40828
rect 12213 40826 12269 40828
rect 12293 40826 12349 40828
rect 12053 40774 12099 40826
rect 12099 40774 12109 40826
rect 12133 40774 12163 40826
rect 12163 40774 12175 40826
rect 12175 40774 12189 40826
rect 12213 40774 12227 40826
rect 12227 40774 12239 40826
rect 12239 40774 12269 40826
rect 12293 40774 12303 40826
rect 12303 40774 12349 40826
rect 12053 40772 12109 40774
rect 12133 40772 12189 40774
rect 12213 40772 12269 40774
rect 12293 40772 12349 40774
rect 16492 40826 16548 40828
rect 16572 40826 16628 40828
rect 16652 40826 16708 40828
rect 16732 40826 16788 40828
rect 16492 40774 16538 40826
rect 16538 40774 16548 40826
rect 16572 40774 16602 40826
rect 16602 40774 16614 40826
rect 16614 40774 16628 40826
rect 16652 40774 16666 40826
rect 16666 40774 16678 40826
rect 16678 40774 16708 40826
rect 16732 40774 16742 40826
rect 16742 40774 16788 40826
rect 16492 40772 16548 40774
rect 16572 40772 16628 40774
rect 16652 40772 16708 40774
rect 16732 40772 16788 40774
rect 18050 40568 18106 40624
rect 5394 40282 5450 40284
rect 5474 40282 5530 40284
rect 5554 40282 5610 40284
rect 5634 40282 5690 40284
rect 5394 40230 5440 40282
rect 5440 40230 5450 40282
rect 5474 40230 5504 40282
rect 5504 40230 5516 40282
rect 5516 40230 5530 40282
rect 5554 40230 5568 40282
rect 5568 40230 5580 40282
rect 5580 40230 5610 40282
rect 5634 40230 5644 40282
rect 5644 40230 5690 40282
rect 5394 40228 5450 40230
rect 5474 40228 5530 40230
rect 5554 40228 5610 40230
rect 5634 40228 5690 40230
rect 9833 40282 9889 40284
rect 9913 40282 9969 40284
rect 9993 40282 10049 40284
rect 10073 40282 10129 40284
rect 9833 40230 9879 40282
rect 9879 40230 9889 40282
rect 9913 40230 9943 40282
rect 9943 40230 9955 40282
rect 9955 40230 9969 40282
rect 9993 40230 10007 40282
rect 10007 40230 10019 40282
rect 10019 40230 10049 40282
rect 10073 40230 10083 40282
rect 10083 40230 10129 40282
rect 9833 40228 9889 40230
rect 9913 40228 9969 40230
rect 9993 40228 10049 40230
rect 10073 40228 10129 40230
rect 14272 40282 14328 40284
rect 14352 40282 14408 40284
rect 14432 40282 14488 40284
rect 14512 40282 14568 40284
rect 14272 40230 14318 40282
rect 14318 40230 14328 40282
rect 14352 40230 14382 40282
rect 14382 40230 14394 40282
rect 14394 40230 14408 40282
rect 14432 40230 14446 40282
rect 14446 40230 14458 40282
rect 14458 40230 14488 40282
rect 14512 40230 14522 40282
rect 14522 40230 14568 40282
rect 14272 40228 14328 40230
rect 14352 40228 14408 40230
rect 14432 40228 14488 40230
rect 14512 40228 14568 40230
rect 3175 39738 3231 39740
rect 3255 39738 3311 39740
rect 3335 39738 3391 39740
rect 3415 39738 3471 39740
rect 3175 39686 3221 39738
rect 3221 39686 3231 39738
rect 3255 39686 3285 39738
rect 3285 39686 3297 39738
rect 3297 39686 3311 39738
rect 3335 39686 3349 39738
rect 3349 39686 3361 39738
rect 3361 39686 3391 39738
rect 3415 39686 3425 39738
rect 3425 39686 3471 39738
rect 3175 39684 3231 39686
rect 3255 39684 3311 39686
rect 3335 39684 3391 39686
rect 3415 39684 3471 39686
rect 7614 39738 7670 39740
rect 7694 39738 7750 39740
rect 7774 39738 7830 39740
rect 7854 39738 7910 39740
rect 7614 39686 7660 39738
rect 7660 39686 7670 39738
rect 7694 39686 7724 39738
rect 7724 39686 7736 39738
rect 7736 39686 7750 39738
rect 7774 39686 7788 39738
rect 7788 39686 7800 39738
rect 7800 39686 7830 39738
rect 7854 39686 7864 39738
rect 7864 39686 7910 39738
rect 7614 39684 7670 39686
rect 7694 39684 7750 39686
rect 7774 39684 7830 39686
rect 7854 39684 7910 39686
rect 12053 39738 12109 39740
rect 12133 39738 12189 39740
rect 12213 39738 12269 39740
rect 12293 39738 12349 39740
rect 12053 39686 12099 39738
rect 12099 39686 12109 39738
rect 12133 39686 12163 39738
rect 12163 39686 12175 39738
rect 12175 39686 12189 39738
rect 12213 39686 12227 39738
rect 12227 39686 12239 39738
rect 12239 39686 12269 39738
rect 12293 39686 12303 39738
rect 12303 39686 12349 39738
rect 12053 39684 12109 39686
rect 12133 39684 12189 39686
rect 12213 39684 12269 39686
rect 12293 39684 12349 39686
rect 16492 39738 16548 39740
rect 16572 39738 16628 39740
rect 16652 39738 16708 39740
rect 16732 39738 16788 39740
rect 16492 39686 16538 39738
rect 16538 39686 16548 39738
rect 16572 39686 16602 39738
rect 16602 39686 16614 39738
rect 16614 39686 16628 39738
rect 16652 39686 16666 39738
rect 16666 39686 16678 39738
rect 16678 39686 16708 39738
rect 16732 39686 16742 39738
rect 16742 39686 16788 39738
rect 16492 39684 16548 39686
rect 16572 39684 16628 39686
rect 16652 39684 16708 39686
rect 16732 39684 16788 39686
rect 5394 39194 5450 39196
rect 5474 39194 5530 39196
rect 5554 39194 5610 39196
rect 5634 39194 5690 39196
rect 5394 39142 5440 39194
rect 5440 39142 5450 39194
rect 5474 39142 5504 39194
rect 5504 39142 5516 39194
rect 5516 39142 5530 39194
rect 5554 39142 5568 39194
rect 5568 39142 5580 39194
rect 5580 39142 5610 39194
rect 5634 39142 5644 39194
rect 5644 39142 5690 39194
rect 5394 39140 5450 39142
rect 5474 39140 5530 39142
rect 5554 39140 5610 39142
rect 5634 39140 5690 39142
rect 9833 39194 9889 39196
rect 9913 39194 9969 39196
rect 9993 39194 10049 39196
rect 10073 39194 10129 39196
rect 9833 39142 9879 39194
rect 9879 39142 9889 39194
rect 9913 39142 9943 39194
rect 9943 39142 9955 39194
rect 9955 39142 9969 39194
rect 9993 39142 10007 39194
rect 10007 39142 10019 39194
rect 10019 39142 10049 39194
rect 10073 39142 10083 39194
rect 10083 39142 10129 39194
rect 9833 39140 9889 39142
rect 9913 39140 9969 39142
rect 9993 39140 10049 39142
rect 10073 39140 10129 39142
rect 14272 39194 14328 39196
rect 14352 39194 14408 39196
rect 14432 39194 14488 39196
rect 14512 39194 14568 39196
rect 14272 39142 14318 39194
rect 14318 39142 14328 39194
rect 14352 39142 14382 39194
rect 14382 39142 14394 39194
rect 14394 39142 14408 39194
rect 14432 39142 14446 39194
rect 14446 39142 14458 39194
rect 14458 39142 14488 39194
rect 14512 39142 14522 39194
rect 14522 39142 14568 39194
rect 14272 39140 14328 39142
rect 14352 39140 14408 39142
rect 14432 39140 14488 39142
rect 14512 39140 14568 39142
rect 3175 38650 3231 38652
rect 3255 38650 3311 38652
rect 3335 38650 3391 38652
rect 3415 38650 3471 38652
rect 3175 38598 3221 38650
rect 3221 38598 3231 38650
rect 3255 38598 3285 38650
rect 3285 38598 3297 38650
rect 3297 38598 3311 38650
rect 3335 38598 3349 38650
rect 3349 38598 3361 38650
rect 3361 38598 3391 38650
rect 3415 38598 3425 38650
rect 3425 38598 3471 38650
rect 3175 38596 3231 38598
rect 3255 38596 3311 38598
rect 3335 38596 3391 38598
rect 3415 38596 3471 38598
rect 7614 38650 7670 38652
rect 7694 38650 7750 38652
rect 7774 38650 7830 38652
rect 7854 38650 7910 38652
rect 7614 38598 7660 38650
rect 7660 38598 7670 38650
rect 7694 38598 7724 38650
rect 7724 38598 7736 38650
rect 7736 38598 7750 38650
rect 7774 38598 7788 38650
rect 7788 38598 7800 38650
rect 7800 38598 7830 38650
rect 7854 38598 7864 38650
rect 7864 38598 7910 38650
rect 7614 38596 7670 38598
rect 7694 38596 7750 38598
rect 7774 38596 7830 38598
rect 7854 38596 7910 38598
rect 12053 38650 12109 38652
rect 12133 38650 12189 38652
rect 12213 38650 12269 38652
rect 12293 38650 12349 38652
rect 12053 38598 12099 38650
rect 12099 38598 12109 38650
rect 12133 38598 12163 38650
rect 12163 38598 12175 38650
rect 12175 38598 12189 38650
rect 12213 38598 12227 38650
rect 12227 38598 12239 38650
rect 12239 38598 12269 38650
rect 12293 38598 12303 38650
rect 12303 38598 12349 38650
rect 12053 38596 12109 38598
rect 12133 38596 12189 38598
rect 12213 38596 12269 38598
rect 12293 38596 12349 38598
rect 16492 38650 16548 38652
rect 16572 38650 16628 38652
rect 16652 38650 16708 38652
rect 16732 38650 16788 38652
rect 16492 38598 16538 38650
rect 16538 38598 16548 38650
rect 16572 38598 16602 38650
rect 16602 38598 16614 38650
rect 16614 38598 16628 38650
rect 16652 38598 16666 38650
rect 16666 38598 16678 38650
rect 16678 38598 16708 38650
rect 16732 38598 16742 38650
rect 16742 38598 16788 38650
rect 16492 38596 16548 38598
rect 16572 38596 16628 38598
rect 16652 38596 16708 38598
rect 16732 38596 16788 38598
rect 5394 38106 5450 38108
rect 5474 38106 5530 38108
rect 5554 38106 5610 38108
rect 5634 38106 5690 38108
rect 5394 38054 5440 38106
rect 5440 38054 5450 38106
rect 5474 38054 5504 38106
rect 5504 38054 5516 38106
rect 5516 38054 5530 38106
rect 5554 38054 5568 38106
rect 5568 38054 5580 38106
rect 5580 38054 5610 38106
rect 5634 38054 5644 38106
rect 5644 38054 5690 38106
rect 5394 38052 5450 38054
rect 5474 38052 5530 38054
rect 5554 38052 5610 38054
rect 5634 38052 5690 38054
rect 9833 38106 9889 38108
rect 9913 38106 9969 38108
rect 9993 38106 10049 38108
rect 10073 38106 10129 38108
rect 9833 38054 9879 38106
rect 9879 38054 9889 38106
rect 9913 38054 9943 38106
rect 9943 38054 9955 38106
rect 9955 38054 9969 38106
rect 9993 38054 10007 38106
rect 10007 38054 10019 38106
rect 10019 38054 10049 38106
rect 10073 38054 10083 38106
rect 10083 38054 10129 38106
rect 9833 38052 9889 38054
rect 9913 38052 9969 38054
rect 9993 38052 10049 38054
rect 10073 38052 10129 38054
rect 14272 38106 14328 38108
rect 14352 38106 14408 38108
rect 14432 38106 14488 38108
rect 14512 38106 14568 38108
rect 14272 38054 14318 38106
rect 14318 38054 14328 38106
rect 14352 38054 14382 38106
rect 14382 38054 14394 38106
rect 14394 38054 14408 38106
rect 14432 38054 14446 38106
rect 14446 38054 14458 38106
rect 14458 38054 14488 38106
rect 14512 38054 14522 38106
rect 14522 38054 14568 38106
rect 14272 38052 14328 38054
rect 14352 38052 14408 38054
rect 14432 38052 14488 38054
rect 14512 38052 14568 38054
rect 3175 37562 3231 37564
rect 3255 37562 3311 37564
rect 3335 37562 3391 37564
rect 3415 37562 3471 37564
rect 3175 37510 3221 37562
rect 3221 37510 3231 37562
rect 3255 37510 3285 37562
rect 3285 37510 3297 37562
rect 3297 37510 3311 37562
rect 3335 37510 3349 37562
rect 3349 37510 3361 37562
rect 3361 37510 3391 37562
rect 3415 37510 3425 37562
rect 3425 37510 3471 37562
rect 3175 37508 3231 37510
rect 3255 37508 3311 37510
rect 3335 37508 3391 37510
rect 3415 37508 3471 37510
rect 7614 37562 7670 37564
rect 7694 37562 7750 37564
rect 7774 37562 7830 37564
rect 7854 37562 7910 37564
rect 7614 37510 7660 37562
rect 7660 37510 7670 37562
rect 7694 37510 7724 37562
rect 7724 37510 7736 37562
rect 7736 37510 7750 37562
rect 7774 37510 7788 37562
rect 7788 37510 7800 37562
rect 7800 37510 7830 37562
rect 7854 37510 7864 37562
rect 7864 37510 7910 37562
rect 7614 37508 7670 37510
rect 7694 37508 7750 37510
rect 7774 37508 7830 37510
rect 7854 37508 7910 37510
rect 12053 37562 12109 37564
rect 12133 37562 12189 37564
rect 12213 37562 12269 37564
rect 12293 37562 12349 37564
rect 12053 37510 12099 37562
rect 12099 37510 12109 37562
rect 12133 37510 12163 37562
rect 12163 37510 12175 37562
rect 12175 37510 12189 37562
rect 12213 37510 12227 37562
rect 12227 37510 12239 37562
rect 12239 37510 12269 37562
rect 12293 37510 12303 37562
rect 12303 37510 12349 37562
rect 12053 37508 12109 37510
rect 12133 37508 12189 37510
rect 12213 37508 12269 37510
rect 12293 37508 12349 37510
rect 16492 37562 16548 37564
rect 16572 37562 16628 37564
rect 16652 37562 16708 37564
rect 16732 37562 16788 37564
rect 16492 37510 16538 37562
rect 16538 37510 16548 37562
rect 16572 37510 16602 37562
rect 16602 37510 16614 37562
rect 16614 37510 16628 37562
rect 16652 37510 16666 37562
rect 16666 37510 16678 37562
rect 16678 37510 16708 37562
rect 16732 37510 16742 37562
rect 16742 37510 16788 37562
rect 16492 37508 16548 37510
rect 16572 37508 16628 37510
rect 16652 37508 16708 37510
rect 16732 37508 16788 37510
rect 5394 37018 5450 37020
rect 5474 37018 5530 37020
rect 5554 37018 5610 37020
rect 5634 37018 5690 37020
rect 5394 36966 5440 37018
rect 5440 36966 5450 37018
rect 5474 36966 5504 37018
rect 5504 36966 5516 37018
rect 5516 36966 5530 37018
rect 5554 36966 5568 37018
rect 5568 36966 5580 37018
rect 5580 36966 5610 37018
rect 5634 36966 5644 37018
rect 5644 36966 5690 37018
rect 5394 36964 5450 36966
rect 5474 36964 5530 36966
rect 5554 36964 5610 36966
rect 5634 36964 5690 36966
rect 9833 37018 9889 37020
rect 9913 37018 9969 37020
rect 9993 37018 10049 37020
rect 10073 37018 10129 37020
rect 9833 36966 9879 37018
rect 9879 36966 9889 37018
rect 9913 36966 9943 37018
rect 9943 36966 9955 37018
rect 9955 36966 9969 37018
rect 9993 36966 10007 37018
rect 10007 36966 10019 37018
rect 10019 36966 10049 37018
rect 10073 36966 10083 37018
rect 10083 36966 10129 37018
rect 9833 36964 9889 36966
rect 9913 36964 9969 36966
rect 9993 36964 10049 36966
rect 10073 36964 10129 36966
rect 14272 37018 14328 37020
rect 14352 37018 14408 37020
rect 14432 37018 14488 37020
rect 14512 37018 14568 37020
rect 14272 36966 14318 37018
rect 14318 36966 14328 37018
rect 14352 36966 14382 37018
rect 14382 36966 14394 37018
rect 14394 36966 14408 37018
rect 14432 36966 14446 37018
rect 14446 36966 14458 37018
rect 14458 36966 14488 37018
rect 14512 36966 14522 37018
rect 14522 36966 14568 37018
rect 14272 36964 14328 36966
rect 14352 36964 14408 36966
rect 14432 36964 14488 36966
rect 14512 36964 14568 36966
rect 3175 36474 3231 36476
rect 3255 36474 3311 36476
rect 3335 36474 3391 36476
rect 3415 36474 3471 36476
rect 3175 36422 3221 36474
rect 3221 36422 3231 36474
rect 3255 36422 3285 36474
rect 3285 36422 3297 36474
rect 3297 36422 3311 36474
rect 3335 36422 3349 36474
rect 3349 36422 3361 36474
rect 3361 36422 3391 36474
rect 3415 36422 3425 36474
rect 3425 36422 3471 36474
rect 3175 36420 3231 36422
rect 3255 36420 3311 36422
rect 3335 36420 3391 36422
rect 3415 36420 3471 36422
rect 7614 36474 7670 36476
rect 7694 36474 7750 36476
rect 7774 36474 7830 36476
rect 7854 36474 7910 36476
rect 7614 36422 7660 36474
rect 7660 36422 7670 36474
rect 7694 36422 7724 36474
rect 7724 36422 7736 36474
rect 7736 36422 7750 36474
rect 7774 36422 7788 36474
rect 7788 36422 7800 36474
rect 7800 36422 7830 36474
rect 7854 36422 7864 36474
rect 7864 36422 7910 36474
rect 7614 36420 7670 36422
rect 7694 36420 7750 36422
rect 7774 36420 7830 36422
rect 7854 36420 7910 36422
rect 12053 36474 12109 36476
rect 12133 36474 12189 36476
rect 12213 36474 12269 36476
rect 12293 36474 12349 36476
rect 12053 36422 12099 36474
rect 12099 36422 12109 36474
rect 12133 36422 12163 36474
rect 12163 36422 12175 36474
rect 12175 36422 12189 36474
rect 12213 36422 12227 36474
rect 12227 36422 12239 36474
rect 12239 36422 12269 36474
rect 12293 36422 12303 36474
rect 12303 36422 12349 36474
rect 12053 36420 12109 36422
rect 12133 36420 12189 36422
rect 12213 36420 12269 36422
rect 12293 36420 12349 36422
rect 16492 36474 16548 36476
rect 16572 36474 16628 36476
rect 16652 36474 16708 36476
rect 16732 36474 16788 36476
rect 16492 36422 16538 36474
rect 16538 36422 16548 36474
rect 16572 36422 16602 36474
rect 16602 36422 16614 36474
rect 16614 36422 16628 36474
rect 16652 36422 16666 36474
rect 16666 36422 16678 36474
rect 16678 36422 16708 36474
rect 16732 36422 16742 36474
rect 16742 36422 16788 36474
rect 16492 36420 16548 36422
rect 16572 36420 16628 36422
rect 16652 36420 16708 36422
rect 16732 36420 16788 36422
rect 5394 35930 5450 35932
rect 5474 35930 5530 35932
rect 5554 35930 5610 35932
rect 5634 35930 5690 35932
rect 5394 35878 5440 35930
rect 5440 35878 5450 35930
rect 5474 35878 5504 35930
rect 5504 35878 5516 35930
rect 5516 35878 5530 35930
rect 5554 35878 5568 35930
rect 5568 35878 5580 35930
rect 5580 35878 5610 35930
rect 5634 35878 5644 35930
rect 5644 35878 5690 35930
rect 5394 35876 5450 35878
rect 5474 35876 5530 35878
rect 5554 35876 5610 35878
rect 5634 35876 5690 35878
rect 9833 35930 9889 35932
rect 9913 35930 9969 35932
rect 9993 35930 10049 35932
rect 10073 35930 10129 35932
rect 9833 35878 9879 35930
rect 9879 35878 9889 35930
rect 9913 35878 9943 35930
rect 9943 35878 9955 35930
rect 9955 35878 9969 35930
rect 9993 35878 10007 35930
rect 10007 35878 10019 35930
rect 10019 35878 10049 35930
rect 10073 35878 10083 35930
rect 10083 35878 10129 35930
rect 9833 35876 9889 35878
rect 9913 35876 9969 35878
rect 9993 35876 10049 35878
rect 10073 35876 10129 35878
rect 14272 35930 14328 35932
rect 14352 35930 14408 35932
rect 14432 35930 14488 35932
rect 14512 35930 14568 35932
rect 14272 35878 14318 35930
rect 14318 35878 14328 35930
rect 14352 35878 14382 35930
rect 14382 35878 14394 35930
rect 14394 35878 14408 35930
rect 14432 35878 14446 35930
rect 14446 35878 14458 35930
rect 14458 35878 14488 35930
rect 14512 35878 14522 35930
rect 14522 35878 14568 35930
rect 14272 35876 14328 35878
rect 14352 35876 14408 35878
rect 14432 35876 14488 35878
rect 14512 35876 14568 35878
rect 3175 35386 3231 35388
rect 3255 35386 3311 35388
rect 3335 35386 3391 35388
rect 3415 35386 3471 35388
rect 3175 35334 3221 35386
rect 3221 35334 3231 35386
rect 3255 35334 3285 35386
rect 3285 35334 3297 35386
rect 3297 35334 3311 35386
rect 3335 35334 3349 35386
rect 3349 35334 3361 35386
rect 3361 35334 3391 35386
rect 3415 35334 3425 35386
rect 3425 35334 3471 35386
rect 3175 35332 3231 35334
rect 3255 35332 3311 35334
rect 3335 35332 3391 35334
rect 3415 35332 3471 35334
rect 7614 35386 7670 35388
rect 7694 35386 7750 35388
rect 7774 35386 7830 35388
rect 7854 35386 7910 35388
rect 7614 35334 7660 35386
rect 7660 35334 7670 35386
rect 7694 35334 7724 35386
rect 7724 35334 7736 35386
rect 7736 35334 7750 35386
rect 7774 35334 7788 35386
rect 7788 35334 7800 35386
rect 7800 35334 7830 35386
rect 7854 35334 7864 35386
rect 7864 35334 7910 35386
rect 7614 35332 7670 35334
rect 7694 35332 7750 35334
rect 7774 35332 7830 35334
rect 7854 35332 7910 35334
rect 12053 35386 12109 35388
rect 12133 35386 12189 35388
rect 12213 35386 12269 35388
rect 12293 35386 12349 35388
rect 12053 35334 12099 35386
rect 12099 35334 12109 35386
rect 12133 35334 12163 35386
rect 12163 35334 12175 35386
rect 12175 35334 12189 35386
rect 12213 35334 12227 35386
rect 12227 35334 12239 35386
rect 12239 35334 12269 35386
rect 12293 35334 12303 35386
rect 12303 35334 12349 35386
rect 12053 35332 12109 35334
rect 12133 35332 12189 35334
rect 12213 35332 12269 35334
rect 12293 35332 12349 35334
rect 16492 35386 16548 35388
rect 16572 35386 16628 35388
rect 16652 35386 16708 35388
rect 16732 35386 16788 35388
rect 16492 35334 16538 35386
rect 16538 35334 16548 35386
rect 16572 35334 16602 35386
rect 16602 35334 16614 35386
rect 16614 35334 16628 35386
rect 16652 35334 16666 35386
rect 16666 35334 16678 35386
rect 16678 35334 16708 35386
rect 16732 35334 16742 35386
rect 16742 35334 16788 35386
rect 16492 35332 16548 35334
rect 16572 35332 16628 35334
rect 16652 35332 16708 35334
rect 16732 35332 16788 35334
rect 5394 34842 5450 34844
rect 5474 34842 5530 34844
rect 5554 34842 5610 34844
rect 5634 34842 5690 34844
rect 5394 34790 5440 34842
rect 5440 34790 5450 34842
rect 5474 34790 5504 34842
rect 5504 34790 5516 34842
rect 5516 34790 5530 34842
rect 5554 34790 5568 34842
rect 5568 34790 5580 34842
rect 5580 34790 5610 34842
rect 5634 34790 5644 34842
rect 5644 34790 5690 34842
rect 5394 34788 5450 34790
rect 5474 34788 5530 34790
rect 5554 34788 5610 34790
rect 5634 34788 5690 34790
rect 9833 34842 9889 34844
rect 9913 34842 9969 34844
rect 9993 34842 10049 34844
rect 10073 34842 10129 34844
rect 9833 34790 9879 34842
rect 9879 34790 9889 34842
rect 9913 34790 9943 34842
rect 9943 34790 9955 34842
rect 9955 34790 9969 34842
rect 9993 34790 10007 34842
rect 10007 34790 10019 34842
rect 10019 34790 10049 34842
rect 10073 34790 10083 34842
rect 10083 34790 10129 34842
rect 9833 34788 9889 34790
rect 9913 34788 9969 34790
rect 9993 34788 10049 34790
rect 10073 34788 10129 34790
rect 14272 34842 14328 34844
rect 14352 34842 14408 34844
rect 14432 34842 14488 34844
rect 14512 34842 14568 34844
rect 14272 34790 14318 34842
rect 14318 34790 14328 34842
rect 14352 34790 14382 34842
rect 14382 34790 14394 34842
rect 14394 34790 14408 34842
rect 14432 34790 14446 34842
rect 14446 34790 14458 34842
rect 14458 34790 14488 34842
rect 14512 34790 14522 34842
rect 14522 34790 14568 34842
rect 14272 34788 14328 34790
rect 14352 34788 14408 34790
rect 14432 34788 14488 34790
rect 14512 34788 14568 34790
rect 3175 34298 3231 34300
rect 3255 34298 3311 34300
rect 3335 34298 3391 34300
rect 3415 34298 3471 34300
rect 3175 34246 3221 34298
rect 3221 34246 3231 34298
rect 3255 34246 3285 34298
rect 3285 34246 3297 34298
rect 3297 34246 3311 34298
rect 3335 34246 3349 34298
rect 3349 34246 3361 34298
rect 3361 34246 3391 34298
rect 3415 34246 3425 34298
rect 3425 34246 3471 34298
rect 3175 34244 3231 34246
rect 3255 34244 3311 34246
rect 3335 34244 3391 34246
rect 3415 34244 3471 34246
rect 7614 34298 7670 34300
rect 7694 34298 7750 34300
rect 7774 34298 7830 34300
rect 7854 34298 7910 34300
rect 7614 34246 7660 34298
rect 7660 34246 7670 34298
rect 7694 34246 7724 34298
rect 7724 34246 7736 34298
rect 7736 34246 7750 34298
rect 7774 34246 7788 34298
rect 7788 34246 7800 34298
rect 7800 34246 7830 34298
rect 7854 34246 7864 34298
rect 7864 34246 7910 34298
rect 7614 34244 7670 34246
rect 7694 34244 7750 34246
rect 7774 34244 7830 34246
rect 7854 34244 7910 34246
rect 12053 34298 12109 34300
rect 12133 34298 12189 34300
rect 12213 34298 12269 34300
rect 12293 34298 12349 34300
rect 12053 34246 12099 34298
rect 12099 34246 12109 34298
rect 12133 34246 12163 34298
rect 12163 34246 12175 34298
rect 12175 34246 12189 34298
rect 12213 34246 12227 34298
rect 12227 34246 12239 34298
rect 12239 34246 12269 34298
rect 12293 34246 12303 34298
rect 12303 34246 12349 34298
rect 12053 34244 12109 34246
rect 12133 34244 12189 34246
rect 12213 34244 12269 34246
rect 12293 34244 12349 34246
rect 16492 34298 16548 34300
rect 16572 34298 16628 34300
rect 16652 34298 16708 34300
rect 16732 34298 16788 34300
rect 16492 34246 16538 34298
rect 16538 34246 16548 34298
rect 16572 34246 16602 34298
rect 16602 34246 16614 34298
rect 16614 34246 16628 34298
rect 16652 34246 16666 34298
rect 16666 34246 16678 34298
rect 16678 34246 16708 34298
rect 16732 34246 16742 34298
rect 16742 34246 16788 34298
rect 16492 34244 16548 34246
rect 16572 34244 16628 34246
rect 16652 34244 16708 34246
rect 16732 34244 16788 34246
rect 5394 33754 5450 33756
rect 5474 33754 5530 33756
rect 5554 33754 5610 33756
rect 5634 33754 5690 33756
rect 5394 33702 5440 33754
rect 5440 33702 5450 33754
rect 5474 33702 5504 33754
rect 5504 33702 5516 33754
rect 5516 33702 5530 33754
rect 5554 33702 5568 33754
rect 5568 33702 5580 33754
rect 5580 33702 5610 33754
rect 5634 33702 5644 33754
rect 5644 33702 5690 33754
rect 5394 33700 5450 33702
rect 5474 33700 5530 33702
rect 5554 33700 5610 33702
rect 5634 33700 5690 33702
rect 9833 33754 9889 33756
rect 9913 33754 9969 33756
rect 9993 33754 10049 33756
rect 10073 33754 10129 33756
rect 9833 33702 9879 33754
rect 9879 33702 9889 33754
rect 9913 33702 9943 33754
rect 9943 33702 9955 33754
rect 9955 33702 9969 33754
rect 9993 33702 10007 33754
rect 10007 33702 10019 33754
rect 10019 33702 10049 33754
rect 10073 33702 10083 33754
rect 10083 33702 10129 33754
rect 9833 33700 9889 33702
rect 9913 33700 9969 33702
rect 9993 33700 10049 33702
rect 10073 33700 10129 33702
rect 14272 33754 14328 33756
rect 14352 33754 14408 33756
rect 14432 33754 14488 33756
rect 14512 33754 14568 33756
rect 14272 33702 14318 33754
rect 14318 33702 14328 33754
rect 14352 33702 14382 33754
rect 14382 33702 14394 33754
rect 14394 33702 14408 33754
rect 14432 33702 14446 33754
rect 14446 33702 14458 33754
rect 14458 33702 14488 33754
rect 14512 33702 14522 33754
rect 14522 33702 14568 33754
rect 14272 33700 14328 33702
rect 14352 33700 14408 33702
rect 14432 33700 14488 33702
rect 14512 33700 14568 33702
rect 3175 33210 3231 33212
rect 3255 33210 3311 33212
rect 3335 33210 3391 33212
rect 3415 33210 3471 33212
rect 3175 33158 3221 33210
rect 3221 33158 3231 33210
rect 3255 33158 3285 33210
rect 3285 33158 3297 33210
rect 3297 33158 3311 33210
rect 3335 33158 3349 33210
rect 3349 33158 3361 33210
rect 3361 33158 3391 33210
rect 3415 33158 3425 33210
rect 3425 33158 3471 33210
rect 3175 33156 3231 33158
rect 3255 33156 3311 33158
rect 3335 33156 3391 33158
rect 3415 33156 3471 33158
rect 7614 33210 7670 33212
rect 7694 33210 7750 33212
rect 7774 33210 7830 33212
rect 7854 33210 7910 33212
rect 7614 33158 7660 33210
rect 7660 33158 7670 33210
rect 7694 33158 7724 33210
rect 7724 33158 7736 33210
rect 7736 33158 7750 33210
rect 7774 33158 7788 33210
rect 7788 33158 7800 33210
rect 7800 33158 7830 33210
rect 7854 33158 7864 33210
rect 7864 33158 7910 33210
rect 7614 33156 7670 33158
rect 7694 33156 7750 33158
rect 7774 33156 7830 33158
rect 7854 33156 7910 33158
rect 12053 33210 12109 33212
rect 12133 33210 12189 33212
rect 12213 33210 12269 33212
rect 12293 33210 12349 33212
rect 12053 33158 12099 33210
rect 12099 33158 12109 33210
rect 12133 33158 12163 33210
rect 12163 33158 12175 33210
rect 12175 33158 12189 33210
rect 12213 33158 12227 33210
rect 12227 33158 12239 33210
rect 12239 33158 12269 33210
rect 12293 33158 12303 33210
rect 12303 33158 12349 33210
rect 12053 33156 12109 33158
rect 12133 33156 12189 33158
rect 12213 33156 12269 33158
rect 12293 33156 12349 33158
rect 16492 33210 16548 33212
rect 16572 33210 16628 33212
rect 16652 33210 16708 33212
rect 16732 33210 16788 33212
rect 16492 33158 16538 33210
rect 16538 33158 16548 33210
rect 16572 33158 16602 33210
rect 16602 33158 16614 33210
rect 16614 33158 16628 33210
rect 16652 33158 16666 33210
rect 16666 33158 16678 33210
rect 16678 33158 16708 33210
rect 16732 33158 16742 33210
rect 16742 33158 16788 33210
rect 16492 33156 16548 33158
rect 16572 33156 16628 33158
rect 16652 33156 16708 33158
rect 16732 33156 16788 33158
rect 5394 32666 5450 32668
rect 5474 32666 5530 32668
rect 5554 32666 5610 32668
rect 5634 32666 5690 32668
rect 5394 32614 5440 32666
rect 5440 32614 5450 32666
rect 5474 32614 5504 32666
rect 5504 32614 5516 32666
rect 5516 32614 5530 32666
rect 5554 32614 5568 32666
rect 5568 32614 5580 32666
rect 5580 32614 5610 32666
rect 5634 32614 5644 32666
rect 5644 32614 5690 32666
rect 5394 32612 5450 32614
rect 5474 32612 5530 32614
rect 5554 32612 5610 32614
rect 5634 32612 5690 32614
rect 9833 32666 9889 32668
rect 9913 32666 9969 32668
rect 9993 32666 10049 32668
rect 10073 32666 10129 32668
rect 9833 32614 9879 32666
rect 9879 32614 9889 32666
rect 9913 32614 9943 32666
rect 9943 32614 9955 32666
rect 9955 32614 9969 32666
rect 9993 32614 10007 32666
rect 10007 32614 10019 32666
rect 10019 32614 10049 32666
rect 10073 32614 10083 32666
rect 10083 32614 10129 32666
rect 9833 32612 9889 32614
rect 9913 32612 9969 32614
rect 9993 32612 10049 32614
rect 10073 32612 10129 32614
rect 14272 32666 14328 32668
rect 14352 32666 14408 32668
rect 14432 32666 14488 32668
rect 14512 32666 14568 32668
rect 14272 32614 14318 32666
rect 14318 32614 14328 32666
rect 14352 32614 14382 32666
rect 14382 32614 14394 32666
rect 14394 32614 14408 32666
rect 14432 32614 14446 32666
rect 14446 32614 14458 32666
rect 14458 32614 14488 32666
rect 14512 32614 14522 32666
rect 14522 32614 14568 32666
rect 14272 32612 14328 32614
rect 14352 32612 14408 32614
rect 14432 32612 14488 32614
rect 14512 32612 14568 32614
rect 3175 32122 3231 32124
rect 3255 32122 3311 32124
rect 3335 32122 3391 32124
rect 3415 32122 3471 32124
rect 3175 32070 3221 32122
rect 3221 32070 3231 32122
rect 3255 32070 3285 32122
rect 3285 32070 3297 32122
rect 3297 32070 3311 32122
rect 3335 32070 3349 32122
rect 3349 32070 3361 32122
rect 3361 32070 3391 32122
rect 3415 32070 3425 32122
rect 3425 32070 3471 32122
rect 3175 32068 3231 32070
rect 3255 32068 3311 32070
rect 3335 32068 3391 32070
rect 3415 32068 3471 32070
rect 7614 32122 7670 32124
rect 7694 32122 7750 32124
rect 7774 32122 7830 32124
rect 7854 32122 7910 32124
rect 7614 32070 7660 32122
rect 7660 32070 7670 32122
rect 7694 32070 7724 32122
rect 7724 32070 7736 32122
rect 7736 32070 7750 32122
rect 7774 32070 7788 32122
rect 7788 32070 7800 32122
rect 7800 32070 7830 32122
rect 7854 32070 7864 32122
rect 7864 32070 7910 32122
rect 7614 32068 7670 32070
rect 7694 32068 7750 32070
rect 7774 32068 7830 32070
rect 7854 32068 7910 32070
rect 12053 32122 12109 32124
rect 12133 32122 12189 32124
rect 12213 32122 12269 32124
rect 12293 32122 12349 32124
rect 12053 32070 12099 32122
rect 12099 32070 12109 32122
rect 12133 32070 12163 32122
rect 12163 32070 12175 32122
rect 12175 32070 12189 32122
rect 12213 32070 12227 32122
rect 12227 32070 12239 32122
rect 12239 32070 12269 32122
rect 12293 32070 12303 32122
rect 12303 32070 12349 32122
rect 12053 32068 12109 32070
rect 12133 32068 12189 32070
rect 12213 32068 12269 32070
rect 12293 32068 12349 32070
rect 16492 32122 16548 32124
rect 16572 32122 16628 32124
rect 16652 32122 16708 32124
rect 16732 32122 16788 32124
rect 16492 32070 16538 32122
rect 16538 32070 16548 32122
rect 16572 32070 16602 32122
rect 16602 32070 16614 32122
rect 16614 32070 16628 32122
rect 16652 32070 16666 32122
rect 16666 32070 16678 32122
rect 16678 32070 16708 32122
rect 16732 32070 16742 32122
rect 16742 32070 16788 32122
rect 16492 32068 16548 32070
rect 16572 32068 16628 32070
rect 16652 32068 16708 32070
rect 16732 32068 16788 32070
rect 5394 31578 5450 31580
rect 5474 31578 5530 31580
rect 5554 31578 5610 31580
rect 5634 31578 5690 31580
rect 5394 31526 5440 31578
rect 5440 31526 5450 31578
rect 5474 31526 5504 31578
rect 5504 31526 5516 31578
rect 5516 31526 5530 31578
rect 5554 31526 5568 31578
rect 5568 31526 5580 31578
rect 5580 31526 5610 31578
rect 5634 31526 5644 31578
rect 5644 31526 5690 31578
rect 5394 31524 5450 31526
rect 5474 31524 5530 31526
rect 5554 31524 5610 31526
rect 5634 31524 5690 31526
rect 9833 31578 9889 31580
rect 9913 31578 9969 31580
rect 9993 31578 10049 31580
rect 10073 31578 10129 31580
rect 9833 31526 9879 31578
rect 9879 31526 9889 31578
rect 9913 31526 9943 31578
rect 9943 31526 9955 31578
rect 9955 31526 9969 31578
rect 9993 31526 10007 31578
rect 10007 31526 10019 31578
rect 10019 31526 10049 31578
rect 10073 31526 10083 31578
rect 10083 31526 10129 31578
rect 9833 31524 9889 31526
rect 9913 31524 9969 31526
rect 9993 31524 10049 31526
rect 10073 31524 10129 31526
rect 14272 31578 14328 31580
rect 14352 31578 14408 31580
rect 14432 31578 14488 31580
rect 14512 31578 14568 31580
rect 14272 31526 14318 31578
rect 14318 31526 14328 31578
rect 14352 31526 14382 31578
rect 14382 31526 14394 31578
rect 14394 31526 14408 31578
rect 14432 31526 14446 31578
rect 14446 31526 14458 31578
rect 14458 31526 14488 31578
rect 14512 31526 14522 31578
rect 14522 31526 14568 31578
rect 14272 31524 14328 31526
rect 14352 31524 14408 31526
rect 14432 31524 14488 31526
rect 14512 31524 14568 31526
rect 3175 31034 3231 31036
rect 3255 31034 3311 31036
rect 3335 31034 3391 31036
rect 3415 31034 3471 31036
rect 3175 30982 3221 31034
rect 3221 30982 3231 31034
rect 3255 30982 3285 31034
rect 3285 30982 3297 31034
rect 3297 30982 3311 31034
rect 3335 30982 3349 31034
rect 3349 30982 3361 31034
rect 3361 30982 3391 31034
rect 3415 30982 3425 31034
rect 3425 30982 3471 31034
rect 3175 30980 3231 30982
rect 3255 30980 3311 30982
rect 3335 30980 3391 30982
rect 3415 30980 3471 30982
rect 7614 31034 7670 31036
rect 7694 31034 7750 31036
rect 7774 31034 7830 31036
rect 7854 31034 7910 31036
rect 7614 30982 7660 31034
rect 7660 30982 7670 31034
rect 7694 30982 7724 31034
rect 7724 30982 7736 31034
rect 7736 30982 7750 31034
rect 7774 30982 7788 31034
rect 7788 30982 7800 31034
rect 7800 30982 7830 31034
rect 7854 30982 7864 31034
rect 7864 30982 7910 31034
rect 7614 30980 7670 30982
rect 7694 30980 7750 30982
rect 7774 30980 7830 30982
rect 7854 30980 7910 30982
rect 12053 31034 12109 31036
rect 12133 31034 12189 31036
rect 12213 31034 12269 31036
rect 12293 31034 12349 31036
rect 12053 30982 12099 31034
rect 12099 30982 12109 31034
rect 12133 30982 12163 31034
rect 12163 30982 12175 31034
rect 12175 30982 12189 31034
rect 12213 30982 12227 31034
rect 12227 30982 12239 31034
rect 12239 30982 12269 31034
rect 12293 30982 12303 31034
rect 12303 30982 12349 31034
rect 12053 30980 12109 30982
rect 12133 30980 12189 30982
rect 12213 30980 12269 30982
rect 12293 30980 12349 30982
rect 16492 31034 16548 31036
rect 16572 31034 16628 31036
rect 16652 31034 16708 31036
rect 16732 31034 16788 31036
rect 16492 30982 16538 31034
rect 16538 30982 16548 31034
rect 16572 30982 16602 31034
rect 16602 30982 16614 31034
rect 16614 30982 16628 31034
rect 16652 30982 16666 31034
rect 16666 30982 16678 31034
rect 16678 30982 16708 31034
rect 16732 30982 16742 31034
rect 16742 30982 16788 31034
rect 16492 30980 16548 30982
rect 16572 30980 16628 30982
rect 16652 30980 16708 30982
rect 16732 30980 16788 30982
rect 5394 30490 5450 30492
rect 5474 30490 5530 30492
rect 5554 30490 5610 30492
rect 5634 30490 5690 30492
rect 5394 30438 5440 30490
rect 5440 30438 5450 30490
rect 5474 30438 5504 30490
rect 5504 30438 5516 30490
rect 5516 30438 5530 30490
rect 5554 30438 5568 30490
rect 5568 30438 5580 30490
rect 5580 30438 5610 30490
rect 5634 30438 5644 30490
rect 5644 30438 5690 30490
rect 5394 30436 5450 30438
rect 5474 30436 5530 30438
rect 5554 30436 5610 30438
rect 5634 30436 5690 30438
rect 9833 30490 9889 30492
rect 9913 30490 9969 30492
rect 9993 30490 10049 30492
rect 10073 30490 10129 30492
rect 9833 30438 9879 30490
rect 9879 30438 9889 30490
rect 9913 30438 9943 30490
rect 9943 30438 9955 30490
rect 9955 30438 9969 30490
rect 9993 30438 10007 30490
rect 10007 30438 10019 30490
rect 10019 30438 10049 30490
rect 10073 30438 10083 30490
rect 10083 30438 10129 30490
rect 9833 30436 9889 30438
rect 9913 30436 9969 30438
rect 9993 30436 10049 30438
rect 10073 30436 10129 30438
rect 14272 30490 14328 30492
rect 14352 30490 14408 30492
rect 14432 30490 14488 30492
rect 14512 30490 14568 30492
rect 14272 30438 14318 30490
rect 14318 30438 14328 30490
rect 14352 30438 14382 30490
rect 14382 30438 14394 30490
rect 14394 30438 14408 30490
rect 14432 30438 14446 30490
rect 14446 30438 14458 30490
rect 14458 30438 14488 30490
rect 14512 30438 14522 30490
rect 14522 30438 14568 30490
rect 14272 30436 14328 30438
rect 14352 30436 14408 30438
rect 14432 30436 14488 30438
rect 14512 30436 14568 30438
rect 3175 29946 3231 29948
rect 3255 29946 3311 29948
rect 3335 29946 3391 29948
rect 3415 29946 3471 29948
rect 3175 29894 3221 29946
rect 3221 29894 3231 29946
rect 3255 29894 3285 29946
rect 3285 29894 3297 29946
rect 3297 29894 3311 29946
rect 3335 29894 3349 29946
rect 3349 29894 3361 29946
rect 3361 29894 3391 29946
rect 3415 29894 3425 29946
rect 3425 29894 3471 29946
rect 3175 29892 3231 29894
rect 3255 29892 3311 29894
rect 3335 29892 3391 29894
rect 3415 29892 3471 29894
rect 7614 29946 7670 29948
rect 7694 29946 7750 29948
rect 7774 29946 7830 29948
rect 7854 29946 7910 29948
rect 7614 29894 7660 29946
rect 7660 29894 7670 29946
rect 7694 29894 7724 29946
rect 7724 29894 7736 29946
rect 7736 29894 7750 29946
rect 7774 29894 7788 29946
rect 7788 29894 7800 29946
rect 7800 29894 7830 29946
rect 7854 29894 7864 29946
rect 7864 29894 7910 29946
rect 7614 29892 7670 29894
rect 7694 29892 7750 29894
rect 7774 29892 7830 29894
rect 7854 29892 7910 29894
rect 12053 29946 12109 29948
rect 12133 29946 12189 29948
rect 12213 29946 12269 29948
rect 12293 29946 12349 29948
rect 12053 29894 12099 29946
rect 12099 29894 12109 29946
rect 12133 29894 12163 29946
rect 12163 29894 12175 29946
rect 12175 29894 12189 29946
rect 12213 29894 12227 29946
rect 12227 29894 12239 29946
rect 12239 29894 12269 29946
rect 12293 29894 12303 29946
rect 12303 29894 12349 29946
rect 12053 29892 12109 29894
rect 12133 29892 12189 29894
rect 12213 29892 12269 29894
rect 12293 29892 12349 29894
rect 16492 29946 16548 29948
rect 16572 29946 16628 29948
rect 16652 29946 16708 29948
rect 16732 29946 16788 29948
rect 16492 29894 16538 29946
rect 16538 29894 16548 29946
rect 16572 29894 16602 29946
rect 16602 29894 16614 29946
rect 16614 29894 16628 29946
rect 16652 29894 16666 29946
rect 16666 29894 16678 29946
rect 16678 29894 16708 29946
rect 16732 29894 16742 29946
rect 16742 29894 16788 29946
rect 16492 29892 16548 29894
rect 16572 29892 16628 29894
rect 16652 29892 16708 29894
rect 16732 29892 16788 29894
rect 5394 29402 5450 29404
rect 5474 29402 5530 29404
rect 5554 29402 5610 29404
rect 5634 29402 5690 29404
rect 5394 29350 5440 29402
rect 5440 29350 5450 29402
rect 5474 29350 5504 29402
rect 5504 29350 5516 29402
rect 5516 29350 5530 29402
rect 5554 29350 5568 29402
rect 5568 29350 5580 29402
rect 5580 29350 5610 29402
rect 5634 29350 5644 29402
rect 5644 29350 5690 29402
rect 5394 29348 5450 29350
rect 5474 29348 5530 29350
rect 5554 29348 5610 29350
rect 5634 29348 5690 29350
rect 9833 29402 9889 29404
rect 9913 29402 9969 29404
rect 9993 29402 10049 29404
rect 10073 29402 10129 29404
rect 9833 29350 9879 29402
rect 9879 29350 9889 29402
rect 9913 29350 9943 29402
rect 9943 29350 9955 29402
rect 9955 29350 9969 29402
rect 9993 29350 10007 29402
rect 10007 29350 10019 29402
rect 10019 29350 10049 29402
rect 10073 29350 10083 29402
rect 10083 29350 10129 29402
rect 9833 29348 9889 29350
rect 9913 29348 9969 29350
rect 9993 29348 10049 29350
rect 10073 29348 10129 29350
rect 14272 29402 14328 29404
rect 14352 29402 14408 29404
rect 14432 29402 14488 29404
rect 14512 29402 14568 29404
rect 14272 29350 14318 29402
rect 14318 29350 14328 29402
rect 14352 29350 14382 29402
rect 14382 29350 14394 29402
rect 14394 29350 14408 29402
rect 14432 29350 14446 29402
rect 14446 29350 14458 29402
rect 14458 29350 14488 29402
rect 14512 29350 14522 29402
rect 14522 29350 14568 29402
rect 14272 29348 14328 29350
rect 14352 29348 14408 29350
rect 14432 29348 14488 29350
rect 14512 29348 14568 29350
rect 3175 28858 3231 28860
rect 3255 28858 3311 28860
rect 3335 28858 3391 28860
rect 3415 28858 3471 28860
rect 3175 28806 3221 28858
rect 3221 28806 3231 28858
rect 3255 28806 3285 28858
rect 3285 28806 3297 28858
rect 3297 28806 3311 28858
rect 3335 28806 3349 28858
rect 3349 28806 3361 28858
rect 3361 28806 3391 28858
rect 3415 28806 3425 28858
rect 3425 28806 3471 28858
rect 3175 28804 3231 28806
rect 3255 28804 3311 28806
rect 3335 28804 3391 28806
rect 3415 28804 3471 28806
rect 7614 28858 7670 28860
rect 7694 28858 7750 28860
rect 7774 28858 7830 28860
rect 7854 28858 7910 28860
rect 7614 28806 7660 28858
rect 7660 28806 7670 28858
rect 7694 28806 7724 28858
rect 7724 28806 7736 28858
rect 7736 28806 7750 28858
rect 7774 28806 7788 28858
rect 7788 28806 7800 28858
rect 7800 28806 7830 28858
rect 7854 28806 7864 28858
rect 7864 28806 7910 28858
rect 7614 28804 7670 28806
rect 7694 28804 7750 28806
rect 7774 28804 7830 28806
rect 7854 28804 7910 28806
rect 12053 28858 12109 28860
rect 12133 28858 12189 28860
rect 12213 28858 12269 28860
rect 12293 28858 12349 28860
rect 12053 28806 12099 28858
rect 12099 28806 12109 28858
rect 12133 28806 12163 28858
rect 12163 28806 12175 28858
rect 12175 28806 12189 28858
rect 12213 28806 12227 28858
rect 12227 28806 12239 28858
rect 12239 28806 12269 28858
rect 12293 28806 12303 28858
rect 12303 28806 12349 28858
rect 12053 28804 12109 28806
rect 12133 28804 12189 28806
rect 12213 28804 12269 28806
rect 12293 28804 12349 28806
rect 16492 28858 16548 28860
rect 16572 28858 16628 28860
rect 16652 28858 16708 28860
rect 16732 28858 16788 28860
rect 16492 28806 16538 28858
rect 16538 28806 16548 28858
rect 16572 28806 16602 28858
rect 16602 28806 16614 28858
rect 16614 28806 16628 28858
rect 16652 28806 16666 28858
rect 16666 28806 16678 28858
rect 16678 28806 16708 28858
rect 16732 28806 16742 28858
rect 16742 28806 16788 28858
rect 16492 28804 16548 28806
rect 16572 28804 16628 28806
rect 16652 28804 16708 28806
rect 16732 28804 16788 28806
rect 5394 28314 5450 28316
rect 5474 28314 5530 28316
rect 5554 28314 5610 28316
rect 5634 28314 5690 28316
rect 5394 28262 5440 28314
rect 5440 28262 5450 28314
rect 5474 28262 5504 28314
rect 5504 28262 5516 28314
rect 5516 28262 5530 28314
rect 5554 28262 5568 28314
rect 5568 28262 5580 28314
rect 5580 28262 5610 28314
rect 5634 28262 5644 28314
rect 5644 28262 5690 28314
rect 5394 28260 5450 28262
rect 5474 28260 5530 28262
rect 5554 28260 5610 28262
rect 5634 28260 5690 28262
rect 9833 28314 9889 28316
rect 9913 28314 9969 28316
rect 9993 28314 10049 28316
rect 10073 28314 10129 28316
rect 9833 28262 9879 28314
rect 9879 28262 9889 28314
rect 9913 28262 9943 28314
rect 9943 28262 9955 28314
rect 9955 28262 9969 28314
rect 9993 28262 10007 28314
rect 10007 28262 10019 28314
rect 10019 28262 10049 28314
rect 10073 28262 10083 28314
rect 10083 28262 10129 28314
rect 9833 28260 9889 28262
rect 9913 28260 9969 28262
rect 9993 28260 10049 28262
rect 10073 28260 10129 28262
rect 14272 28314 14328 28316
rect 14352 28314 14408 28316
rect 14432 28314 14488 28316
rect 14512 28314 14568 28316
rect 14272 28262 14318 28314
rect 14318 28262 14328 28314
rect 14352 28262 14382 28314
rect 14382 28262 14394 28314
rect 14394 28262 14408 28314
rect 14432 28262 14446 28314
rect 14446 28262 14458 28314
rect 14458 28262 14488 28314
rect 14512 28262 14522 28314
rect 14522 28262 14568 28314
rect 14272 28260 14328 28262
rect 14352 28260 14408 28262
rect 14432 28260 14488 28262
rect 14512 28260 14568 28262
rect 3175 27770 3231 27772
rect 3255 27770 3311 27772
rect 3335 27770 3391 27772
rect 3415 27770 3471 27772
rect 3175 27718 3221 27770
rect 3221 27718 3231 27770
rect 3255 27718 3285 27770
rect 3285 27718 3297 27770
rect 3297 27718 3311 27770
rect 3335 27718 3349 27770
rect 3349 27718 3361 27770
rect 3361 27718 3391 27770
rect 3415 27718 3425 27770
rect 3425 27718 3471 27770
rect 3175 27716 3231 27718
rect 3255 27716 3311 27718
rect 3335 27716 3391 27718
rect 3415 27716 3471 27718
rect 7614 27770 7670 27772
rect 7694 27770 7750 27772
rect 7774 27770 7830 27772
rect 7854 27770 7910 27772
rect 7614 27718 7660 27770
rect 7660 27718 7670 27770
rect 7694 27718 7724 27770
rect 7724 27718 7736 27770
rect 7736 27718 7750 27770
rect 7774 27718 7788 27770
rect 7788 27718 7800 27770
rect 7800 27718 7830 27770
rect 7854 27718 7864 27770
rect 7864 27718 7910 27770
rect 7614 27716 7670 27718
rect 7694 27716 7750 27718
rect 7774 27716 7830 27718
rect 7854 27716 7910 27718
rect 12053 27770 12109 27772
rect 12133 27770 12189 27772
rect 12213 27770 12269 27772
rect 12293 27770 12349 27772
rect 12053 27718 12099 27770
rect 12099 27718 12109 27770
rect 12133 27718 12163 27770
rect 12163 27718 12175 27770
rect 12175 27718 12189 27770
rect 12213 27718 12227 27770
rect 12227 27718 12239 27770
rect 12239 27718 12269 27770
rect 12293 27718 12303 27770
rect 12303 27718 12349 27770
rect 12053 27716 12109 27718
rect 12133 27716 12189 27718
rect 12213 27716 12269 27718
rect 12293 27716 12349 27718
rect 16492 27770 16548 27772
rect 16572 27770 16628 27772
rect 16652 27770 16708 27772
rect 16732 27770 16788 27772
rect 16492 27718 16538 27770
rect 16538 27718 16548 27770
rect 16572 27718 16602 27770
rect 16602 27718 16614 27770
rect 16614 27718 16628 27770
rect 16652 27718 16666 27770
rect 16666 27718 16678 27770
rect 16678 27718 16708 27770
rect 16732 27718 16742 27770
rect 16742 27718 16788 27770
rect 16492 27716 16548 27718
rect 16572 27716 16628 27718
rect 16652 27716 16708 27718
rect 16732 27716 16788 27718
rect 5394 27226 5450 27228
rect 5474 27226 5530 27228
rect 5554 27226 5610 27228
rect 5634 27226 5690 27228
rect 5394 27174 5440 27226
rect 5440 27174 5450 27226
rect 5474 27174 5504 27226
rect 5504 27174 5516 27226
rect 5516 27174 5530 27226
rect 5554 27174 5568 27226
rect 5568 27174 5580 27226
rect 5580 27174 5610 27226
rect 5634 27174 5644 27226
rect 5644 27174 5690 27226
rect 5394 27172 5450 27174
rect 5474 27172 5530 27174
rect 5554 27172 5610 27174
rect 5634 27172 5690 27174
rect 9833 27226 9889 27228
rect 9913 27226 9969 27228
rect 9993 27226 10049 27228
rect 10073 27226 10129 27228
rect 9833 27174 9879 27226
rect 9879 27174 9889 27226
rect 9913 27174 9943 27226
rect 9943 27174 9955 27226
rect 9955 27174 9969 27226
rect 9993 27174 10007 27226
rect 10007 27174 10019 27226
rect 10019 27174 10049 27226
rect 10073 27174 10083 27226
rect 10083 27174 10129 27226
rect 9833 27172 9889 27174
rect 9913 27172 9969 27174
rect 9993 27172 10049 27174
rect 10073 27172 10129 27174
rect 14272 27226 14328 27228
rect 14352 27226 14408 27228
rect 14432 27226 14488 27228
rect 14512 27226 14568 27228
rect 14272 27174 14318 27226
rect 14318 27174 14328 27226
rect 14352 27174 14382 27226
rect 14382 27174 14394 27226
rect 14394 27174 14408 27226
rect 14432 27174 14446 27226
rect 14446 27174 14458 27226
rect 14458 27174 14488 27226
rect 14512 27174 14522 27226
rect 14522 27174 14568 27226
rect 14272 27172 14328 27174
rect 14352 27172 14408 27174
rect 14432 27172 14488 27174
rect 14512 27172 14568 27174
rect 3175 26682 3231 26684
rect 3255 26682 3311 26684
rect 3335 26682 3391 26684
rect 3415 26682 3471 26684
rect 3175 26630 3221 26682
rect 3221 26630 3231 26682
rect 3255 26630 3285 26682
rect 3285 26630 3297 26682
rect 3297 26630 3311 26682
rect 3335 26630 3349 26682
rect 3349 26630 3361 26682
rect 3361 26630 3391 26682
rect 3415 26630 3425 26682
rect 3425 26630 3471 26682
rect 3175 26628 3231 26630
rect 3255 26628 3311 26630
rect 3335 26628 3391 26630
rect 3415 26628 3471 26630
rect 7614 26682 7670 26684
rect 7694 26682 7750 26684
rect 7774 26682 7830 26684
rect 7854 26682 7910 26684
rect 7614 26630 7660 26682
rect 7660 26630 7670 26682
rect 7694 26630 7724 26682
rect 7724 26630 7736 26682
rect 7736 26630 7750 26682
rect 7774 26630 7788 26682
rect 7788 26630 7800 26682
rect 7800 26630 7830 26682
rect 7854 26630 7864 26682
rect 7864 26630 7910 26682
rect 7614 26628 7670 26630
rect 7694 26628 7750 26630
rect 7774 26628 7830 26630
rect 7854 26628 7910 26630
rect 12053 26682 12109 26684
rect 12133 26682 12189 26684
rect 12213 26682 12269 26684
rect 12293 26682 12349 26684
rect 12053 26630 12099 26682
rect 12099 26630 12109 26682
rect 12133 26630 12163 26682
rect 12163 26630 12175 26682
rect 12175 26630 12189 26682
rect 12213 26630 12227 26682
rect 12227 26630 12239 26682
rect 12239 26630 12269 26682
rect 12293 26630 12303 26682
rect 12303 26630 12349 26682
rect 12053 26628 12109 26630
rect 12133 26628 12189 26630
rect 12213 26628 12269 26630
rect 12293 26628 12349 26630
rect 16492 26682 16548 26684
rect 16572 26682 16628 26684
rect 16652 26682 16708 26684
rect 16732 26682 16788 26684
rect 16492 26630 16538 26682
rect 16538 26630 16548 26682
rect 16572 26630 16602 26682
rect 16602 26630 16614 26682
rect 16614 26630 16628 26682
rect 16652 26630 16666 26682
rect 16666 26630 16678 26682
rect 16678 26630 16708 26682
rect 16732 26630 16742 26682
rect 16742 26630 16788 26682
rect 16492 26628 16548 26630
rect 16572 26628 16628 26630
rect 16652 26628 16708 26630
rect 16732 26628 16788 26630
rect 5394 26138 5450 26140
rect 5474 26138 5530 26140
rect 5554 26138 5610 26140
rect 5634 26138 5690 26140
rect 5394 26086 5440 26138
rect 5440 26086 5450 26138
rect 5474 26086 5504 26138
rect 5504 26086 5516 26138
rect 5516 26086 5530 26138
rect 5554 26086 5568 26138
rect 5568 26086 5580 26138
rect 5580 26086 5610 26138
rect 5634 26086 5644 26138
rect 5644 26086 5690 26138
rect 5394 26084 5450 26086
rect 5474 26084 5530 26086
rect 5554 26084 5610 26086
rect 5634 26084 5690 26086
rect 9833 26138 9889 26140
rect 9913 26138 9969 26140
rect 9993 26138 10049 26140
rect 10073 26138 10129 26140
rect 9833 26086 9879 26138
rect 9879 26086 9889 26138
rect 9913 26086 9943 26138
rect 9943 26086 9955 26138
rect 9955 26086 9969 26138
rect 9993 26086 10007 26138
rect 10007 26086 10019 26138
rect 10019 26086 10049 26138
rect 10073 26086 10083 26138
rect 10083 26086 10129 26138
rect 9833 26084 9889 26086
rect 9913 26084 9969 26086
rect 9993 26084 10049 26086
rect 10073 26084 10129 26086
rect 14272 26138 14328 26140
rect 14352 26138 14408 26140
rect 14432 26138 14488 26140
rect 14512 26138 14568 26140
rect 14272 26086 14318 26138
rect 14318 26086 14328 26138
rect 14352 26086 14382 26138
rect 14382 26086 14394 26138
rect 14394 26086 14408 26138
rect 14432 26086 14446 26138
rect 14446 26086 14458 26138
rect 14458 26086 14488 26138
rect 14512 26086 14522 26138
rect 14522 26086 14568 26138
rect 14272 26084 14328 26086
rect 14352 26084 14408 26086
rect 14432 26084 14488 26086
rect 14512 26084 14568 26086
rect 3175 25594 3231 25596
rect 3255 25594 3311 25596
rect 3335 25594 3391 25596
rect 3415 25594 3471 25596
rect 3175 25542 3221 25594
rect 3221 25542 3231 25594
rect 3255 25542 3285 25594
rect 3285 25542 3297 25594
rect 3297 25542 3311 25594
rect 3335 25542 3349 25594
rect 3349 25542 3361 25594
rect 3361 25542 3391 25594
rect 3415 25542 3425 25594
rect 3425 25542 3471 25594
rect 3175 25540 3231 25542
rect 3255 25540 3311 25542
rect 3335 25540 3391 25542
rect 3415 25540 3471 25542
rect 7614 25594 7670 25596
rect 7694 25594 7750 25596
rect 7774 25594 7830 25596
rect 7854 25594 7910 25596
rect 7614 25542 7660 25594
rect 7660 25542 7670 25594
rect 7694 25542 7724 25594
rect 7724 25542 7736 25594
rect 7736 25542 7750 25594
rect 7774 25542 7788 25594
rect 7788 25542 7800 25594
rect 7800 25542 7830 25594
rect 7854 25542 7864 25594
rect 7864 25542 7910 25594
rect 7614 25540 7670 25542
rect 7694 25540 7750 25542
rect 7774 25540 7830 25542
rect 7854 25540 7910 25542
rect 12053 25594 12109 25596
rect 12133 25594 12189 25596
rect 12213 25594 12269 25596
rect 12293 25594 12349 25596
rect 12053 25542 12099 25594
rect 12099 25542 12109 25594
rect 12133 25542 12163 25594
rect 12163 25542 12175 25594
rect 12175 25542 12189 25594
rect 12213 25542 12227 25594
rect 12227 25542 12239 25594
rect 12239 25542 12269 25594
rect 12293 25542 12303 25594
rect 12303 25542 12349 25594
rect 12053 25540 12109 25542
rect 12133 25540 12189 25542
rect 12213 25540 12269 25542
rect 12293 25540 12349 25542
rect 16492 25594 16548 25596
rect 16572 25594 16628 25596
rect 16652 25594 16708 25596
rect 16732 25594 16788 25596
rect 16492 25542 16538 25594
rect 16538 25542 16548 25594
rect 16572 25542 16602 25594
rect 16602 25542 16614 25594
rect 16614 25542 16628 25594
rect 16652 25542 16666 25594
rect 16666 25542 16678 25594
rect 16678 25542 16708 25594
rect 16732 25542 16742 25594
rect 16742 25542 16788 25594
rect 16492 25540 16548 25542
rect 16572 25540 16628 25542
rect 16652 25540 16708 25542
rect 16732 25540 16788 25542
rect 5394 25050 5450 25052
rect 5474 25050 5530 25052
rect 5554 25050 5610 25052
rect 5634 25050 5690 25052
rect 5394 24998 5440 25050
rect 5440 24998 5450 25050
rect 5474 24998 5504 25050
rect 5504 24998 5516 25050
rect 5516 24998 5530 25050
rect 5554 24998 5568 25050
rect 5568 24998 5580 25050
rect 5580 24998 5610 25050
rect 5634 24998 5644 25050
rect 5644 24998 5690 25050
rect 5394 24996 5450 24998
rect 5474 24996 5530 24998
rect 5554 24996 5610 24998
rect 5634 24996 5690 24998
rect 9833 25050 9889 25052
rect 9913 25050 9969 25052
rect 9993 25050 10049 25052
rect 10073 25050 10129 25052
rect 9833 24998 9879 25050
rect 9879 24998 9889 25050
rect 9913 24998 9943 25050
rect 9943 24998 9955 25050
rect 9955 24998 9969 25050
rect 9993 24998 10007 25050
rect 10007 24998 10019 25050
rect 10019 24998 10049 25050
rect 10073 24998 10083 25050
rect 10083 24998 10129 25050
rect 9833 24996 9889 24998
rect 9913 24996 9969 24998
rect 9993 24996 10049 24998
rect 10073 24996 10129 24998
rect 14272 25050 14328 25052
rect 14352 25050 14408 25052
rect 14432 25050 14488 25052
rect 14512 25050 14568 25052
rect 14272 24998 14318 25050
rect 14318 24998 14328 25050
rect 14352 24998 14382 25050
rect 14382 24998 14394 25050
rect 14394 24998 14408 25050
rect 14432 24998 14446 25050
rect 14446 24998 14458 25050
rect 14458 24998 14488 25050
rect 14512 24998 14522 25050
rect 14522 24998 14568 25050
rect 14272 24996 14328 24998
rect 14352 24996 14408 24998
rect 14432 24996 14488 24998
rect 14512 24996 14568 24998
rect 3175 24506 3231 24508
rect 3255 24506 3311 24508
rect 3335 24506 3391 24508
rect 3415 24506 3471 24508
rect 3175 24454 3221 24506
rect 3221 24454 3231 24506
rect 3255 24454 3285 24506
rect 3285 24454 3297 24506
rect 3297 24454 3311 24506
rect 3335 24454 3349 24506
rect 3349 24454 3361 24506
rect 3361 24454 3391 24506
rect 3415 24454 3425 24506
rect 3425 24454 3471 24506
rect 3175 24452 3231 24454
rect 3255 24452 3311 24454
rect 3335 24452 3391 24454
rect 3415 24452 3471 24454
rect 7614 24506 7670 24508
rect 7694 24506 7750 24508
rect 7774 24506 7830 24508
rect 7854 24506 7910 24508
rect 7614 24454 7660 24506
rect 7660 24454 7670 24506
rect 7694 24454 7724 24506
rect 7724 24454 7736 24506
rect 7736 24454 7750 24506
rect 7774 24454 7788 24506
rect 7788 24454 7800 24506
rect 7800 24454 7830 24506
rect 7854 24454 7864 24506
rect 7864 24454 7910 24506
rect 7614 24452 7670 24454
rect 7694 24452 7750 24454
rect 7774 24452 7830 24454
rect 7854 24452 7910 24454
rect 12053 24506 12109 24508
rect 12133 24506 12189 24508
rect 12213 24506 12269 24508
rect 12293 24506 12349 24508
rect 12053 24454 12099 24506
rect 12099 24454 12109 24506
rect 12133 24454 12163 24506
rect 12163 24454 12175 24506
rect 12175 24454 12189 24506
rect 12213 24454 12227 24506
rect 12227 24454 12239 24506
rect 12239 24454 12269 24506
rect 12293 24454 12303 24506
rect 12303 24454 12349 24506
rect 12053 24452 12109 24454
rect 12133 24452 12189 24454
rect 12213 24452 12269 24454
rect 12293 24452 12349 24454
rect 16492 24506 16548 24508
rect 16572 24506 16628 24508
rect 16652 24506 16708 24508
rect 16732 24506 16788 24508
rect 16492 24454 16538 24506
rect 16538 24454 16548 24506
rect 16572 24454 16602 24506
rect 16602 24454 16614 24506
rect 16614 24454 16628 24506
rect 16652 24454 16666 24506
rect 16666 24454 16678 24506
rect 16678 24454 16708 24506
rect 16732 24454 16742 24506
rect 16742 24454 16788 24506
rect 16492 24452 16548 24454
rect 16572 24452 16628 24454
rect 16652 24452 16708 24454
rect 16732 24452 16788 24454
rect 5394 23962 5450 23964
rect 5474 23962 5530 23964
rect 5554 23962 5610 23964
rect 5634 23962 5690 23964
rect 5394 23910 5440 23962
rect 5440 23910 5450 23962
rect 5474 23910 5504 23962
rect 5504 23910 5516 23962
rect 5516 23910 5530 23962
rect 5554 23910 5568 23962
rect 5568 23910 5580 23962
rect 5580 23910 5610 23962
rect 5634 23910 5644 23962
rect 5644 23910 5690 23962
rect 5394 23908 5450 23910
rect 5474 23908 5530 23910
rect 5554 23908 5610 23910
rect 5634 23908 5690 23910
rect 9833 23962 9889 23964
rect 9913 23962 9969 23964
rect 9993 23962 10049 23964
rect 10073 23962 10129 23964
rect 9833 23910 9879 23962
rect 9879 23910 9889 23962
rect 9913 23910 9943 23962
rect 9943 23910 9955 23962
rect 9955 23910 9969 23962
rect 9993 23910 10007 23962
rect 10007 23910 10019 23962
rect 10019 23910 10049 23962
rect 10073 23910 10083 23962
rect 10083 23910 10129 23962
rect 9833 23908 9889 23910
rect 9913 23908 9969 23910
rect 9993 23908 10049 23910
rect 10073 23908 10129 23910
rect 14272 23962 14328 23964
rect 14352 23962 14408 23964
rect 14432 23962 14488 23964
rect 14512 23962 14568 23964
rect 14272 23910 14318 23962
rect 14318 23910 14328 23962
rect 14352 23910 14382 23962
rect 14382 23910 14394 23962
rect 14394 23910 14408 23962
rect 14432 23910 14446 23962
rect 14446 23910 14458 23962
rect 14458 23910 14488 23962
rect 14512 23910 14522 23962
rect 14522 23910 14568 23962
rect 14272 23908 14328 23910
rect 14352 23908 14408 23910
rect 14432 23908 14488 23910
rect 14512 23908 14568 23910
rect 3175 23418 3231 23420
rect 3255 23418 3311 23420
rect 3335 23418 3391 23420
rect 3415 23418 3471 23420
rect 3175 23366 3221 23418
rect 3221 23366 3231 23418
rect 3255 23366 3285 23418
rect 3285 23366 3297 23418
rect 3297 23366 3311 23418
rect 3335 23366 3349 23418
rect 3349 23366 3361 23418
rect 3361 23366 3391 23418
rect 3415 23366 3425 23418
rect 3425 23366 3471 23418
rect 3175 23364 3231 23366
rect 3255 23364 3311 23366
rect 3335 23364 3391 23366
rect 3415 23364 3471 23366
rect 7614 23418 7670 23420
rect 7694 23418 7750 23420
rect 7774 23418 7830 23420
rect 7854 23418 7910 23420
rect 7614 23366 7660 23418
rect 7660 23366 7670 23418
rect 7694 23366 7724 23418
rect 7724 23366 7736 23418
rect 7736 23366 7750 23418
rect 7774 23366 7788 23418
rect 7788 23366 7800 23418
rect 7800 23366 7830 23418
rect 7854 23366 7864 23418
rect 7864 23366 7910 23418
rect 7614 23364 7670 23366
rect 7694 23364 7750 23366
rect 7774 23364 7830 23366
rect 7854 23364 7910 23366
rect 12053 23418 12109 23420
rect 12133 23418 12189 23420
rect 12213 23418 12269 23420
rect 12293 23418 12349 23420
rect 12053 23366 12099 23418
rect 12099 23366 12109 23418
rect 12133 23366 12163 23418
rect 12163 23366 12175 23418
rect 12175 23366 12189 23418
rect 12213 23366 12227 23418
rect 12227 23366 12239 23418
rect 12239 23366 12269 23418
rect 12293 23366 12303 23418
rect 12303 23366 12349 23418
rect 12053 23364 12109 23366
rect 12133 23364 12189 23366
rect 12213 23364 12269 23366
rect 12293 23364 12349 23366
rect 16492 23418 16548 23420
rect 16572 23418 16628 23420
rect 16652 23418 16708 23420
rect 16732 23418 16788 23420
rect 16492 23366 16538 23418
rect 16538 23366 16548 23418
rect 16572 23366 16602 23418
rect 16602 23366 16614 23418
rect 16614 23366 16628 23418
rect 16652 23366 16666 23418
rect 16666 23366 16678 23418
rect 16678 23366 16708 23418
rect 16732 23366 16742 23418
rect 16742 23366 16788 23418
rect 16492 23364 16548 23366
rect 16572 23364 16628 23366
rect 16652 23364 16708 23366
rect 16732 23364 16788 23366
rect 5394 22874 5450 22876
rect 5474 22874 5530 22876
rect 5554 22874 5610 22876
rect 5634 22874 5690 22876
rect 5394 22822 5440 22874
rect 5440 22822 5450 22874
rect 5474 22822 5504 22874
rect 5504 22822 5516 22874
rect 5516 22822 5530 22874
rect 5554 22822 5568 22874
rect 5568 22822 5580 22874
rect 5580 22822 5610 22874
rect 5634 22822 5644 22874
rect 5644 22822 5690 22874
rect 5394 22820 5450 22822
rect 5474 22820 5530 22822
rect 5554 22820 5610 22822
rect 5634 22820 5690 22822
rect 9833 22874 9889 22876
rect 9913 22874 9969 22876
rect 9993 22874 10049 22876
rect 10073 22874 10129 22876
rect 9833 22822 9879 22874
rect 9879 22822 9889 22874
rect 9913 22822 9943 22874
rect 9943 22822 9955 22874
rect 9955 22822 9969 22874
rect 9993 22822 10007 22874
rect 10007 22822 10019 22874
rect 10019 22822 10049 22874
rect 10073 22822 10083 22874
rect 10083 22822 10129 22874
rect 9833 22820 9889 22822
rect 9913 22820 9969 22822
rect 9993 22820 10049 22822
rect 10073 22820 10129 22822
rect 14272 22874 14328 22876
rect 14352 22874 14408 22876
rect 14432 22874 14488 22876
rect 14512 22874 14568 22876
rect 14272 22822 14318 22874
rect 14318 22822 14328 22874
rect 14352 22822 14382 22874
rect 14382 22822 14394 22874
rect 14394 22822 14408 22874
rect 14432 22822 14446 22874
rect 14446 22822 14458 22874
rect 14458 22822 14488 22874
rect 14512 22822 14522 22874
rect 14522 22822 14568 22874
rect 14272 22820 14328 22822
rect 14352 22820 14408 22822
rect 14432 22820 14488 22822
rect 14512 22820 14568 22822
rect 3175 22330 3231 22332
rect 3255 22330 3311 22332
rect 3335 22330 3391 22332
rect 3415 22330 3471 22332
rect 3175 22278 3221 22330
rect 3221 22278 3231 22330
rect 3255 22278 3285 22330
rect 3285 22278 3297 22330
rect 3297 22278 3311 22330
rect 3335 22278 3349 22330
rect 3349 22278 3361 22330
rect 3361 22278 3391 22330
rect 3415 22278 3425 22330
rect 3425 22278 3471 22330
rect 3175 22276 3231 22278
rect 3255 22276 3311 22278
rect 3335 22276 3391 22278
rect 3415 22276 3471 22278
rect 7614 22330 7670 22332
rect 7694 22330 7750 22332
rect 7774 22330 7830 22332
rect 7854 22330 7910 22332
rect 7614 22278 7660 22330
rect 7660 22278 7670 22330
rect 7694 22278 7724 22330
rect 7724 22278 7736 22330
rect 7736 22278 7750 22330
rect 7774 22278 7788 22330
rect 7788 22278 7800 22330
rect 7800 22278 7830 22330
rect 7854 22278 7864 22330
rect 7864 22278 7910 22330
rect 7614 22276 7670 22278
rect 7694 22276 7750 22278
rect 7774 22276 7830 22278
rect 7854 22276 7910 22278
rect 12053 22330 12109 22332
rect 12133 22330 12189 22332
rect 12213 22330 12269 22332
rect 12293 22330 12349 22332
rect 12053 22278 12099 22330
rect 12099 22278 12109 22330
rect 12133 22278 12163 22330
rect 12163 22278 12175 22330
rect 12175 22278 12189 22330
rect 12213 22278 12227 22330
rect 12227 22278 12239 22330
rect 12239 22278 12269 22330
rect 12293 22278 12303 22330
rect 12303 22278 12349 22330
rect 12053 22276 12109 22278
rect 12133 22276 12189 22278
rect 12213 22276 12269 22278
rect 12293 22276 12349 22278
rect 16492 22330 16548 22332
rect 16572 22330 16628 22332
rect 16652 22330 16708 22332
rect 16732 22330 16788 22332
rect 16492 22278 16538 22330
rect 16538 22278 16548 22330
rect 16572 22278 16602 22330
rect 16602 22278 16614 22330
rect 16614 22278 16628 22330
rect 16652 22278 16666 22330
rect 16666 22278 16678 22330
rect 16678 22278 16708 22330
rect 16732 22278 16742 22330
rect 16742 22278 16788 22330
rect 16492 22276 16548 22278
rect 16572 22276 16628 22278
rect 16652 22276 16708 22278
rect 16732 22276 16788 22278
rect 5394 21786 5450 21788
rect 5474 21786 5530 21788
rect 5554 21786 5610 21788
rect 5634 21786 5690 21788
rect 5394 21734 5440 21786
rect 5440 21734 5450 21786
rect 5474 21734 5504 21786
rect 5504 21734 5516 21786
rect 5516 21734 5530 21786
rect 5554 21734 5568 21786
rect 5568 21734 5580 21786
rect 5580 21734 5610 21786
rect 5634 21734 5644 21786
rect 5644 21734 5690 21786
rect 5394 21732 5450 21734
rect 5474 21732 5530 21734
rect 5554 21732 5610 21734
rect 5634 21732 5690 21734
rect 9833 21786 9889 21788
rect 9913 21786 9969 21788
rect 9993 21786 10049 21788
rect 10073 21786 10129 21788
rect 9833 21734 9879 21786
rect 9879 21734 9889 21786
rect 9913 21734 9943 21786
rect 9943 21734 9955 21786
rect 9955 21734 9969 21786
rect 9993 21734 10007 21786
rect 10007 21734 10019 21786
rect 10019 21734 10049 21786
rect 10073 21734 10083 21786
rect 10083 21734 10129 21786
rect 9833 21732 9889 21734
rect 9913 21732 9969 21734
rect 9993 21732 10049 21734
rect 10073 21732 10129 21734
rect 14272 21786 14328 21788
rect 14352 21786 14408 21788
rect 14432 21786 14488 21788
rect 14512 21786 14568 21788
rect 14272 21734 14318 21786
rect 14318 21734 14328 21786
rect 14352 21734 14382 21786
rect 14382 21734 14394 21786
rect 14394 21734 14408 21786
rect 14432 21734 14446 21786
rect 14446 21734 14458 21786
rect 14458 21734 14488 21786
rect 14512 21734 14522 21786
rect 14522 21734 14568 21786
rect 14272 21732 14328 21734
rect 14352 21732 14408 21734
rect 14432 21732 14488 21734
rect 14512 21732 14568 21734
rect 3175 21242 3231 21244
rect 3255 21242 3311 21244
rect 3335 21242 3391 21244
rect 3415 21242 3471 21244
rect 3175 21190 3221 21242
rect 3221 21190 3231 21242
rect 3255 21190 3285 21242
rect 3285 21190 3297 21242
rect 3297 21190 3311 21242
rect 3335 21190 3349 21242
rect 3349 21190 3361 21242
rect 3361 21190 3391 21242
rect 3415 21190 3425 21242
rect 3425 21190 3471 21242
rect 3175 21188 3231 21190
rect 3255 21188 3311 21190
rect 3335 21188 3391 21190
rect 3415 21188 3471 21190
rect 7614 21242 7670 21244
rect 7694 21242 7750 21244
rect 7774 21242 7830 21244
rect 7854 21242 7910 21244
rect 7614 21190 7660 21242
rect 7660 21190 7670 21242
rect 7694 21190 7724 21242
rect 7724 21190 7736 21242
rect 7736 21190 7750 21242
rect 7774 21190 7788 21242
rect 7788 21190 7800 21242
rect 7800 21190 7830 21242
rect 7854 21190 7864 21242
rect 7864 21190 7910 21242
rect 7614 21188 7670 21190
rect 7694 21188 7750 21190
rect 7774 21188 7830 21190
rect 7854 21188 7910 21190
rect 12053 21242 12109 21244
rect 12133 21242 12189 21244
rect 12213 21242 12269 21244
rect 12293 21242 12349 21244
rect 12053 21190 12099 21242
rect 12099 21190 12109 21242
rect 12133 21190 12163 21242
rect 12163 21190 12175 21242
rect 12175 21190 12189 21242
rect 12213 21190 12227 21242
rect 12227 21190 12239 21242
rect 12239 21190 12269 21242
rect 12293 21190 12303 21242
rect 12303 21190 12349 21242
rect 12053 21188 12109 21190
rect 12133 21188 12189 21190
rect 12213 21188 12269 21190
rect 12293 21188 12349 21190
rect 16492 21242 16548 21244
rect 16572 21242 16628 21244
rect 16652 21242 16708 21244
rect 16732 21242 16788 21244
rect 16492 21190 16538 21242
rect 16538 21190 16548 21242
rect 16572 21190 16602 21242
rect 16602 21190 16614 21242
rect 16614 21190 16628 21242
rect 16652 21190 16666 21242
rect 16666 21190 16678 21242
rect 16678 21190 16708 21242
rect 16732 21190 16742 21242
rect 16742 21190 16788 21242
rect 16492 21188 16548 21190
rect 16572 21188 16628 21190
rect 16652 21188 16708 21190
rect 16732 21188 16788 21190
rect 5394 20698 5450 20700
rect 5474 20698 5530 20700
rect 5554 20698 5610 20700
rect 5634 20698 5690 20700
rect 5394 20646 5440 20698
rect 5440 20646 5450 20698
rect 5474 20646 5504 20698
rect 5504 20646 5516 20698
rect 5516 20646 5530 20698
rect 5554 20646 5568 20698
rect 5568 20646 5580 20698
rect 5580 20646 5610 20698
rect 5634 20646 5644 20698
rect 5644 20646 5690 20698
rect 5394 20644 5450 20646
rect 5474 20644 5530 20646
rect 5554 20644 5610 20646
rect 5634 20644 5690 20646
rect 9833 20698 9889 20700
rect 9913 20698 9969 20700
rect 9993 20698 10049 20700
rect 10073 20698 10129 20700
rect 9833 20646 9879 20698
rect 9879 20646 9889 20698
rect 9913 20646 9943 20698
rect 9943 20646 9955 20698
rect 9955 20646 9969 20698
rect 9993 20646 10007 20698
rect 10007 20646 10019 20698
rect 10019 20646 10049 20698
rect 10073 20646 10083 20698
rect 10083 20646 10129 20698
rect 9833 20644 9889 20646
rect 9913 20644 9969 20646
rect 9993 20644 10049 20646
rect 10073 20644 10129 20646
rect 14272 20698 14328 20700
rect 14352 20698 14408 20700
rect 14432 20698 14488 20700
rect 14512 20698 14568 20700
rect 14272 20646 14318 20698
rect 14318 20646 14328 20698
rect 14352 20646 14382 20698
rect 14382 20646 14394 20698
rect 14394 20646 14408 20698
rect 14432 20646 14446 20698
rect 14446 20646 14458 20698
rect 14458 20646 14488 20698
rect 14512 20646 14522 20698
rect 14522 20646 14568 20698
rect 14272 20644 14328 20646
rect 14352 20644 14408 20646
rect 14432 20644 14488 20646
rect 14512 20644 14568 20646
rect 3175 20154 3231 20156
rect 3255 20154 3311 20156
rect 3335 20154 3391 20156
rect 3415 20154 3471 20156
rect 3175 20102 3221 20154
rect 3221 20102 3231 20154
rect 3255 20102 3285 20154
rect 3285 20102 3297 20154
rect 3297 20102 3311 20154
rect 3335 20102 3349 20154
rect 3349 20102 3361 20154
rect 3361 20102 3391 20154
rect 3415 20102 3425 20154
rect 3425 20102 3471 20154
rect 3175 20100 3231 20102
rect 3255 20100 3311 20102
rect 3335 20100 3391 20102
rect 3415 20100 3471 20102
rect 7614 20154 7670 20156
rect 7694 20154 7750 20156
rect 7774 20154 7830 20156
rect 7854 20154 7910 20156
rect 7614 20102 7660 20154
rect 7660 20102 7670 20154
rect 7694 20102 7724 20154
rect 7724 20102 7736 20154
rect 7736 20102 7750 20154
rect 7774 20102 7788 20154
rect 7788 20102 7800 20154
rect 7800 20102 7830 20154
rect 7854 20102 7864 20154
rect 7864 20102 7910 20154
rect 7614 20100 7670 20102
rect 7694 20100 7750 20102
rect 7774 20100 7830 20102
rect 7854 20100 7910 20102
rect 12053 20154 12109 20156
rect 12133 20154 12189 20156
rect 12213 20154 12269 20156
rect 12293 20154 12349 20156
rect 12053 20102 12099 20154
rect 12099 20102 12109 20154
rect 12133 20102 12163 20154
rect 12163 20102 12175 20154
rect 12175 20102 12189 20154
rect 12213 20102 12227 20154
rect 12227 20102 12239 20154
rect 12239 20102 12269 20154
rect 12293 20102 12303 20154
rect 12303 20102 12349 20154
rect 12053 20100 12109 20102
rect 12133 20100 12189 20102
rect 12213 20100 12269 20102
rect 12293 20100 12349 20102
rect 16492 20154 16548 20156
rect 16572 20154 16628 20156
rect 16652 20154 16708 20156
rect 16732 20154 16788 20156
rect 16492 20102 16538 20154
rect 16538 20102 16548 20154
rect 16572 20102 16602 20154
rect 16602 20102 16614 20154
rect 16614 20102 16628 20154
rect 16652 20102 16666 20154
rect 16666 20102 16678 20154
rect 16678 20102 16708 20154
rect 16732 20102 16742 20154
rect 16742 20102 16788 20154
rect 16492 20100 16548 20102
rect 16572 20100 16628 20102
rect 16652 20100 16708 20102
rect 16732 20100 16788 20102
rect 5394 19610 5450 19612
rect 5474 19610 5530 19612
rect 5554 19610 5610 19612
rect 5634 19610 5690 19612
rect 5394 19558 5440 19610
rect 5440 19558 5450 19610
rect 5474 19558 5504 19610
rect 5504 19558 5516 19610
rect 5516 19558 5530 19610
rect 5554 19558 5568 19610
rect 5568 19558 5580 19610
rect 5580 19558 5610 19610
rect 5634 19558 5644 19610
rect 5644 19558 5690 19610
rect 5394 19556 5450 19558
rect 5474 19556 5530 19558
rect 5554 19556 5610 19558
rect 5634 19556 5690 19558
rect 9833 19610 9889 19612
rect 9913 19610 9969 19612
rect 9993 19610 10049 19612
rect 10073 19610 10129 19612
rect 9833 19558 9879 19610
rect 9879 19558 9889 19610
rect 9913 19558 9943 19610
rect 9943 19558 9955 19610
rect 9955 19558 9969 19610
rect 9993 19558 10007 19610
rect 10007 19558 10019 19610
rect 10019 19558 10049 19610
rect 10073 19558 10083 19610
rect 10083 19558 10129 19610
rect 9833 19556 9889 19558
rect 9913 19556 9969 19558
rect 9993 19556 10049 19558
rect 10073 19556 10129 19558
rect 14272 19610 14328 19612
rect 14352 19610 14408 19612
rect 14432 19610 14488 19612
rect 14512 19610 14568 19612
rect 14272 19558 14318 19610
rect 14318 19558 14328 19610
rect 14352 19558 14382 19610
rect 14382 19558 14394 19610
rect 14394 19558 14408 19610
rect 14432 19558 14446 19610
rect 14446 19558 14458 19610
rect 14458 19558 14488 19610
rect 14512 19558 14522 19610
rect 14522 19558 14568 19610
rect 14272 19556 14328 19558
rect 14352 19556 14408 19558
rect 14432 19556 14488 19558
rect 14512 19556 14568 19558
rect 3175 19066 3231 19068
rect 3255 19066 3311 19068
rect 3335 19066 3391 19068
rect 3415 19066 3471 19068
rect 3175 19014 3221 19066
rect 3221 19014 3231 19066
rect 3255 19014 3285 19066
rect 3285 19014 3297 19066
rect 3297 19014 3311 19066
rect 3335 19014 3349 19066
rect 3349 19014 3361 19066
rect 3361 19014 3391 19066
rect 3415 19014 3425 19066
rect 3425 19014 3471 19066
rect 3175 19012 3231 19014
rect 3255 19012 3311 19014
rect 3335 19012 3391 19014
rect 3415 19012 3471 19014
rect 7614 19066 7670 19068
rect 7694 19066 7750 19068
rect 7774 19066 7830 19068
rect 7854 19066 7910 19068
rect 7614 19014 7660 19066
rect 7660 19014 7670 19066
rect 7694 19014 7724 19066
rect 7724 19014 7736 19066
rect 7736 19014 7750 19066
rect 7774 19014 7788 19066
rect 7788 19014 7800 19066
rect 7800 19014 7830 19066
rect 7854 19014 7864 19066
rect 7864 19014 7910 19066
rect 7614 19012 7670 19014
rect 7694 19012 7750 19014
rect 7774 19012 7830 19014
rect 7854 19012 7910 19014
rect 12053 19066 12109 19068
rect 12133 19066 12189 19068
rect 12213 19066 12269 19068
rect 12293 19066 12349 19068
rect 12053 19014 12099 19066
rect 12099 19014 12109 19066
rect 12133 19014 12163 19066
rect 12163 19014 12175 19066
rect 12175 19014 12189 19066
rect 12213 19014 12227 19066
rect 12227 19014 12239 19066
rect 12239 19014 12269 19066
rect 12293 19014 12303 19066
rect 12303 19014 12349 19066
rect 12053 19012 12109 19014
rect 12133 19012 12189 19014
rect 12213 19012 12269 19014
rect 12293 19012 12349 19014
rect 16492 19066 16548 19068
rect 16572 19066 16628 19068
rect 16652 19066 16708 19068
rect 16732 19066 16788 19068
rect 16492 19014 16538 19066
rect 16538 19014 16548 19066
rect 16572 19014 16602 19066
rect 16602 19014 16614 19066
rect 16614 19014 16628 19066
rect 16652 19014 16666 19066
rect 16666 19014 16678 19066
rect 16678 19014 16708 19066
rect 16732 19014 16742 19066
rect 16742 19014 16788 19066
rect 16492 19012 16548 19014
rect 16572 19012 16628 19014
rect 16652 19012 16708 19014
rect 16732 19012 16788 19014
rect 5394 18522 5450 18524
rect 5474 18522 5530 18524
rect 5554 18522 5610 18524
rect 5634 18522 5690 18524
rect 5394 18470 5440 18522
rect 5440 18470 5450 18522
rect 5474 18470 5504 18522
rect 5504 18470 5516 18522
rect 5516 18470 5530 18522
rect 5554 18470 5568 18522
rect 5568 18470 5580 18522
rect 5580 18470 5610 18522
rect 5634 18470 5644 18522
rect 5644 18470 5690 18522
rect 5394 18468 5450 18470
rect 5474 18468 5530 18470
rect 5554 18468 5610 18470
rect 5634 18468 5690 18470
rect 9833 18522 9889 18524
rect 9913 18522 9969 18524
rect 9993 18522 10049 18524
rect 10073 18522 10129 18524
rect 9833 18470 9879 18522
rect 9879 18470 9889 18522
rect 9913 18470 9943 18522
rect 9943 18470 9955 18522
rect 9955 18470 9969 18522
rect 9993 18470 10007 18522
rect 10007 18470 10019 18522
rect 10019 18470 10049 18522
rect 10073 18470 10083 18522
rect 10083 18470 10129 18522
rect 9833 18468 9889 18470
rect 9913 18468 9969 18470
rect 9993 18468 10049 18470
rect 10073 18468 10129 18470
rect 14272 18522 14328 18524
rect 14352 18522 14408 18524
rect 14432 18522 14488 18524
rect 14512 18522 14568 18524
rect 14272 18470 14318 18522
rect 14318 18470 14328 18522
rect 14352 18470 14382 18522
rect 14382 18470 14394 18522
rect 14394 18470 14408 18522
rect 14432 18470 14446 18522
rect 14446 18470 14458 18522
rect 14458 18470 14488 18522
rect 14512 18470 14522 18522
rect 14522 18470 14568 18522
rect 14272 18468 14328 18470
rect 14352 18468 14408 18470
rect 14432 18468 14488 18470
rect 14512 18468 14568 18470
rect 3175 17978 3231 17980
rect 3255 17978 3311 17980
rect 3335 17978 3391 17980
rect 3415 17978 3471 17980
rect 3175 17926 3221 17978
rect 3221 17926 3231 17978
rect 3255 17926 3285 17978
rect 3285 17926 3297 17978
rect 3297 17926 3311 17978
rect 3335 17926 3349 17978
rect 3349 17926 3361 17978
rect 3361 17926 3391 17978
rect 3415 17926 3425 17978
rect 3425 17926 3471 17978
rect 3175 17924 3231 17926
rect 3255 17924 3311 17926
rect 3335 17924 3391 17926
rect 3415 17924 3471 17926
rect 7614 17978 7670 17980
rect 7694 17978 7750 17980
rect 7774 17978 7830 17980
rect 7854 17978 7910 17980
rect 7614 17926 7660 17978
rect 7660 17926 7670 17978
rect 7694 17926 7724 17978
rect 7724 17926 7736 17978
rect 7736 17926 7750 17978
rect 7774 17926 7788 17978
rect 7788 17926 7800 17978
rect 7800 17926 7830 17978
rect 7854 17926 7864 17978
rect 7864 17926 7910 17978
rect 7614 17924 7670 17926
rect 7694 17924 7750 17926
rect 7774 17924 7830 17926
rect 7854 17924 7910 17926
rect 12053 17978 12109 17980
rect 12133 17978 12189 17980
rect 12213 17978 12269 17980
rect 12293 17978 12349 17980
rect 12053 17926 12099 17978
rect 12099 17926 12109 17978
rect 12133 17926 12163 17978
rect 12163 17926 12175 17978
rect 12175 17926 12189 17978
rect 12213 17926 12227 17978
rect 12227 17926 12239 17978
rect 12239 17926 12269 17978
rect 12293 17926 12303 17978
rect 12303 17926 12349 17978
rect 12053 17924 12109 17926
rect 12133 17924 12189 17926
rect 12213 17924 12269 17926
rect 12293 17924 12349 17926
rect 16492 17978 16548 17980
rect 16572 17978 16628 17980
rect 16652 17978 16708 17980
rect 16732 17978 16788 17980
rect 16492 17926 16538 17978
rect 16538 17926 16548 17978
rect 16572 17926 16602 17978
rect 16602 17926 16614 17978
rect 16614 17926 16628 17978
rect 16652 17926 16666 17978
rect 16666 17926 16678 17978
rect 16678 17926 16708 17978
rect 16732 17926 16742 17978
rect 16742 17926 16788 17978
rect 16492 17924 16548 17926
rect 16572 17924 16628 17926
rect 16652 17924 16708 17926
rect 16732 17924 16788 17926
rect 5394 17434 5450 17436
rect 5474 17434 5530 17436
rect 5554 17434 5610 17436
rect 5634 17434 5690 17436
rect 5394 17382 5440 17434
rect 5440 17382 5450 17434
rect 5474 17382 5504 17434
rect 5504 17382 5516 17434
rect 5516 17382 5530 17434
rect 5554 17382 5568 17434
rect 5568 17382 5580 17434
rect 5580 17382 5610 17434
rect 5634 17382 5644 17434
rect 5644 17382 5690 17434
rect 5394 17380 5450 17382
rect 5474 17380 5530 17382
rect 5554 17380 5610 17382
rect 5634 17380 5690 17382
rect 9833 17434 9889 17436
rect 9913 17434 9969 17436
rect 9993 17434 10049 17436
rect 10073 17434 10129 17436
rect 9833 17382 9879 17434
rect 9879 17382 9889 17434
rect 9913 17382 9943 17434
rect 9943 17382 9955 17434
rect 9955 17382 9969 17434
rect 9993 17382 10007 17434
rect 10007 17382 10019 17434
rect 10019 17382 10049 17434
rect 10073 17382 10083 17434
rect 10083 17382 10129 17434
rect 9833 17380 9889 17382
rect 9913 17380 9969 17382
rect 9993 17380 10049 17382
rect 10073 17380 10129 17382
rect 14272 17434 14328 17436
rect 14352 17434 14408 17436
rect 14432 17434 14488 17436
rect 14512 17434 14568 17436
rect 14272 17382 14318 17434
rect 14318 17382 14328 17434
rect 14352 17382 14382 17434
rect 14382 17382 14394 17434
rect 14394 17382 14408 17434
rect 14432 17382 14446 17434
rect 14446 17382 14458 17434
rect 14458 17382 14488 17434
rect 14512 17382 14522 17434
rect 14522 17382 14568 17434
rect 14272 17380 14328 17382
rect 14352 17380 14408 17382
rect 14432 17380 14488 17382
rect 14512 17380 14568 17382
rect 3175 16890 3231 16892
rect 3255 16890 3311 16892
rect 3335 16890 3391 16892
rect 3415 16890 3471 16892
rect 3175 16838 3221 16890
rect 3221 16838 3231 16890
rect 3255 16838 3285 16890
rect 3285 16838 3297 16890
rect 3297 16838 3311 16890
rect 3335 16838 3349 16890
rect 3349 16838 3361 16890
rect 3361 16838 3391 16890
rect 3415 16838 3425 16890
rect 3425 16838 3471 16890
rect 3175 16836 3231 16838
rect 3255 16836 3311 16838
rect 3335 16836 3391 16838
rect 3415 16836 3471 16838
rect 7614 16890 7670 16892
rect 7694 16890 7750 16892
rect 7774 16890 7830 16892
rect 7854 16890 7910 16892
rect 7614 16838 7660 16890
rect 7660 16838 7670 16890
rect 7694 16838 7724 16890
rect 7724 16838 7736 16890
rect 7736 16838 7750 16890
rect 7774 16838 7788 16890
rect 7788 16838 7800 16890
rect 7800 16838 7830 16890
rect 7854 16838 7864 16890
rect 7864 16838 7910 16890
rect 7614 16836 7670 16838
rect 7694 16836 7750 16838
rect 7774 16836 7830 16838
rect 7854 16836 7910 16838
rect 12053 16890 12109 16892
rect 12133 16890 12189 16892
rect 12213 16890 12269 16892
rect 12293 16890 12349 16892
rect 12053 16838 12099 16890
rect 12099 16838 12109 16890
rect 12133 16838 12163 16890
rect 12163 16838 12175 16890
rect 12175 16838 12189 16890
rect 12213 16838 12227 16890
rect 12227 16838 12239 16890
rect 12239 16838 12269 16890
rect 12293 16838 12303 16890
rect 12303 16838 12349 16890
rect 12053 16836 12109 16838
rect 12133 16836 12189 16838
rect 12213 16836 12269 16838
rect 12293 16836 12349 16838
rect 16492 16890 16548 16892
rect 16572 16890 16628 16892
rect 16652 16890 16708 16892
rect 16732 16890 16788 16892
rect 16492 16838 16538 16890
rect 16538 16838 16548 16890
rect 16572 16838 16602 16890
rect 16602 16838 16614 16890
rect 16614 16838 16628 16890
rect 16652 16838 16666 16890
rect 16666 16838 16678 16890
rect 16678 16838 16708 16890
rect 16732 16838 16742 16890
rect 16742 16838 16788 16890
rect 16492 16836 16548 16838
rect 16572 16836 16628 16838
rect 16652 16836 16708 16838
rect 16732 16836 16788 16838
rect 5394 16346 5450 16348
rect 5474 16346 5530 16348
rect 5554 16346 5610 16348
rect 5634 16346 5690 16348
rect 5394 16294 5440 16346
rect 5440 16294 5450 16346
rect 5474 16294 5504 16346
rect 5504 16294 5516 16346
rect 5516 16294 5530 16346
rect 5554 16294 5568 16346
rect 5568 16294 5580 16346
rect 5580 16294 5610 16346
rect 5634 16294 5644 16346
rect 5644 16294 5690 16346
rect 5394 16292 5450 16294
rect 5474 16292 5530 16294
rect 5554 16292 5610 16294
rect 5634 16292 5690 16294
rect 9833 16346 9889 16348
rect 9913 16346 9969 16348
rect 9993 16346 10049 16348
rect 10073 16346 10129 16348
rect 9833 16294 9879 16346
rect 9879 16294 9889 16346
rect 9913 16294 9943 16346
rect 9943 16294 9955 16346
rect 9955 16294 9969 16346
rect 9993 16294 10007 16346
rect 10007 16294 10019 16346
rect 10019 16294 10049 16346
rect 10073 16294 10083 16346
rect 10083 16294 10129 16346
rect 9833 16292 9889 16294
rect 9913 16292 9969 16294
rect 9993 16292 10049 16294
rect 10073 16292 10129 16294
rect 14272 16346 14328 16348
rect 14352 16346 14408 16348
rect 14432 16346 14488 16348
rect 14512 16346 14568 16348
rect 14272 16294 14318 16346
rect 14318 16294 14328 16346
rect 14352 16294 14382 16346
rect 14382 16294 14394 16346
rect 14394 16294 14408 16346
rect 14432 16294 14446 16346
rect 14446 16294 14458 16346
rect 14458 16294 14488 16346
rect 14512 16294 14522 16346
rect 14522 16294 14568 16346
rect 14272 16292 14328 16294
rect 14352 16292 14408 16294
rect 14432 16292 14488 16294
rect 14512 16292 14568 16294
rect 3175 15802 3231 15804
rect 3255 15802 3311 15804
rect 3335 15802 3391 15804
rect 3415 15802 3471 15804
rect 3175 15750 3221 15802
rect 3221 15750 3231 15802
rect 3255 15750 3285 15802
rect 3285 15750 3297 15802
rect 3297 15750 3311 15802
rect 3335 15750 3349 15802
rect 3349 15750 3361 15802
rect 3361 15750 3391 15802
rect 3415 15750 3425 15802
rect 3425 15750 3471 15802
rect 3175 15748 3231 15750
rect 3255 15748 3311 15750
rect 3335 15748 3391 15750
rect 3415 15748 3471 15750
rect 7614 15802 7670 15804
rect 7694 15802 7750 15804
rect 7774 15802 7830 15804
rect 7854 15802 7910 15804
rect 7614 15750 7660 15802
rect 7660 15750 7670 15802
rect 7694 15750 7724 15802
rect 7724 15750 7736 15802
rect 7736 15750 7750 15802
rect 7774 15750 7788 15802
rect 7788 15750 7800 15802
rect 7800 15750 7830 15802
rect 7854 15750 7864 15802
rect 7864 15750 7910 15802
rect 7614 15748 7670 15750
rect 7694 15748 7750 15750
rect 7774 15748 7830 15750
rect 7854 15748 7910 15750
rect 12053 15802 12109 15804
rect 12133 15802 12189 15804
rect 12213 15802 12269 15804
rect 12293 15802 12349 15804
rect 12053 15750 12099 15802
rect 12099 15750 12109 15802
rect 12133 15750 12163 15802
rect 12163 15750 12175 15802
rect 12175 15750 12189 15802
rect 12213 15750 12227 15802
rect 12227 15750 12239 15802
rect 12239 15750 12269 15802
rect 12293 15750 12303 15802
rect 12303 15750 12349 15802
rect 12053 15748 12109 15750
rect 12133 15748 12189 15750
rect 12213 15748 12269 15750
rect 12293 15748 12349 15750
rect 16492 15802 16548 15804
rect 16572 15802 16628 15804
rect 16652 15802 16708 15804
rect 16732 15802 16788 15804
rect 16492 15750 16538 15802
rect 16538 15750 16548 15802
rect 16572 15750 16602 15802
rect 16602 15750 16614 15802
rect 16614 15750 16628 15802
rect 16652 15750 16666 15802
rect 16666 15750 16678 15802
rect 16678 15750 16708 15802
rect 16732 15750 16742 15802
rect 16742 15750 16788 15802
rect 16492 15748 16548 15750
rect 16572 15748 16628 15750
rect 16652 15748 16708 15750
rect 16732 15748 16788 15750
rect 5394 15258 5450 15260
rect 5474 15258 5530 15260
rect 5554 15258 5610 15260
rect 5634 15258 5690 15260
rect 5394 15206 5440 15258
rect 5440 15206 5450 15258
rect 5474 15206 5504 15258
rect 5504 15206 5516 15258
rect 5516 15206 5530 15258
rect 5554 15206 5568 15258
rect 5568 15206 5580 15258
rect 5580 15206 5610 15258
rect 5634 15206 5644 15258
rect 5644 15206 5690 15258
rect 5394 15204 5450 15206
rect 5474 15204 5530 15206
rect 5554 15204 5610 15206
rect 5634 15204 5690 15206
rect 9833 15258 9889 15260
rect 9913 15258 9969 15260
rect 9993 15258 10049 15260
rect 10073 15258 10129 15260
rect 9833 15206 9879 15258
rect 9879 15206 9889 15258
rect 9913 15206 9943 15258
rect 9943 15206 9955 15258
rect 9955 15206 9969 15258
rect 9993 15206 10007 15258
rect 10007 15206 10019 15258
rect 10019 15206 10049 15258
rect 10073 15206 10083 15258
rect 10083 15206 10129 15258
rect 9833 15204 9889 15206
rect 9913 15204 9969 15206
rect 9993 15204 10049 15206
rect 10073 15204 10129 15206
rect 14272 15258 14328 15260
rect 14352 15258 14408 15260
rect 14432 15258 14488 15260
rect 14512 15258 14568 15260
rect 14272 15206 14318 15258
rect 14318 15206 14328 15258
rect 14352 15206 14382 15258
rect 14382 15206 14394 15258
rect 14394 15206 14408 15258
rect 14432 15206 14446 15258
rect 14446 15206 14458 15258
rect 14458 15206 14488 15258
rect 14512 15206 14522 15258
rect 14522 15206 14568 15258
rect 14272 15204 14328 15206
rect 14352 15204 14408 15206
rect 14432 15204 14488 15206
rect 14512 15204 14568 15206
rect 3175 14714 3231 14716
rect 3255 14714 3311 14716
rect 3335 14714 3391 14716
rect 3415 14714 3471 14716
rect 3175 14662 3221 14714
rect 3221 14662 3231 14714
rect 3255 14662 3285 14714
rect 3285 14662 3297 14714
rect 3297 14662 3311 14714
rect 3335 14662 3349 14714
rect 3349 14662 3361 14714
rect 3361 14662 3391 14714
rect 3415 14662 3425 14714
rect 3425 14662 3471 14714
rect 3175 14660 3231 14662
rect 3255 14660 3311 14662
rect 3335 14660 3391 14662
rect 3415 14660 3471 14662
rect 7614 14714 7670 14716
rect 7694 14714 7750 14716
rect 7774 14714 7830 14716
rect 7854 14714 7910 14716
rect 7614 14662 7660 14714
rect 7660 14662 7670 14714
rect 7694 14662 7724 14714
rect 7724 14662 7736 14714
rect 7736 14662 7750 14714
rect 7774 14662 7788 14714
rect 7788 14662 7800 14714
rect 7800 14662 7830 14714
rect 7854 14662 7864 14714
rect 7864 14662 7910 14714
rect 7614 14660 7670 14662
rect 7694 14660 7750 14662
rect 7774 14660 7830 14662
rect 7854 14660 7910 14662
rect 12053 14714 12109 14716
rect 12133 14714 12189 14716
rect 12213 14714 12269 14716
rect 12293 14714 12349 14716
rect 12053 14662 12099 14714
rect 12099 14662 12109 14714
rect 12133 14662 12163 14714
rect 12163 14662 12175 14714
rect 12175 14662 12189 14714
rect 12213 14662 12227 14714
rect 12227 14662 12239 14714
rect 12239 14662 12269 14714
rect 12293 14662 12303 14714
rect 12303 14662 12349 14714
rect 12053 14660 12109 14662
rect 12133 14660 12189 14662
rect 12213 14660 12269 14662
rect 12293 14660 12349 14662
rect 16492 14714 16548 14716
rect 16572 14714 16628 14716
rect 16652 14714 16708 14716
rect 16732 14714 16788 14716
rect 16492 14662 16538 14714
rect 16538 14662 16548 14714
rect 16572 14662 16602 14714
rect 16602 14662 16614 14714
rect 16614 14662 16628 14714
rect 16652 14662 16666 14714
rect 16666 14662 16678 14714
rect 16678 14662 16708 14714
rect 16732 14662 16742 14714
rect 16742 14662 16788 14714
rect 16492 14660 16548 14662
rect 16572 14660 16628 14662
rect 16652 14660 16708 14662
rect 16732 14660 16788 14662
rect 5394 14170 5450 14172
rect 5474 14170 5530 14172
rect 5554 14170 5610 14172
rect 5634 14170 5690 14172
rect 5394 14118 5440 14170
rect 5440 14118 5450 14170
rect 5474 14118 5504 14170
rect 5504 14118 5516 14170
rect 5516 14118 5530 14170
rect 5554 14118 5568 14170
rect 5568 14118 5580 14170
rect 5580 14118 5610 14170
rect 5634 14118 5644 14170
rect 5644 14118 5690 14170
rect 5394 14116 5450 14118
rect 5474 14116 5530 14118
rect 5554 14116 5610 14118
rect 5634 14116 5690 14118
rect 9833 14170 9889 14172
rect 9913 14170 9969 14172
rect 9993 14170 10049 14172
rect 10073 14170 10129 14172
rect 9833 14118 9879 14170
rect 9879 14118 9889 14170
rect 9913 14118 9943 14170
rect 9943 14118 9955 14170
rect 9955 14118 9969 14170
rect 9993 14118 10007 14170
rect 10007 14118 10019 14170
rect 10019 14118 10049 14170
rect 10073 14118 10083 14170
rect 10083 14118 10129 14170
rect 9833 14116 9889 14118
rect 9913 14116 9969 14118
rect 9993 14116 10049 14118
rect 10073 14116 10129 14118
rect 14272 14170 14328 14172
rect 14352 14170 14408 14172
rect 14432 14170 14488 14172
rect 14512 14170 14568 14172
rect 14272 14118 14318 14170
rect 14318 14118 14328 14170
rect 14352 14118 14382 14170
rect 14382 14118 14394 14170
rect 14394 14118 14408 14170
rect 14432 14118 14446 14170
rect 14446 14118 14458 14170
rect 14458 14118 14488 14170
rect 14512 14118 14522 14170
rect 14522 14118 14568 14170
rect 14272 14116 14328 14118
rect 14352 14116 14408 14118
rect 14432 14116 14488 14118
rect 14512 14116 14568 14118
rect 3175 13626 3231 13628
rect 3255 13626 3311 13628
rect 3335 13626 3391 13628
rect 3415 13626 3471 13628
rect 3175 13574 3221 13626
rect 3221 13574 3231 13626
rect 3255 13574 3285 13626
rect 3285 13574 3297 13626
rect 3297 13574 3311 13626
rect 3335 13574 3349 13626
rect 3349 13574 3361 13626
rect 3361 13574 3391 13626
rect 3415 13574 3425 13626
rect 3425 13574 3471 13626
rect 3175 13572 3231 13574
rect 3255 13572 3311 13574
rect 3335 13572 3391 13574
rect 3415 13572 3471 13574
rect 7614 13626 7670 13628
rect 7694 13626 7750 13628
rect 7774 13626 7830 13628
rect 7854 13626 7910 13628
rect 7614 13574 7660 13626
rect 7660 13574 7670 13626
rect 7694 13574 7724 13626
rect 7724 13574 7736 13626
rect 7736 13574 7750 13626
rect 7774 13574 7788 13626
rect 7788 13574 7800 13626
rect 7800 13574 7830 13626
rect 7854 13574 7864 13626
rect 7864 13574 7910 13626
rect 7614 13572 7670 13574
rect 7694 13572 7750 13574
rect 7774 13572 7830 13574
rect 7854 13572 7910 13574
rect 12053 13626 12109 13628
rect 12133 13626 12189 13628
rect 12213 13626 12269 13628
rect 12293 13626 12349 13628
rect 12053 13574 12099 13626
rect 12099 13574 12109 13626
rect 12133 13574 12163 13626
rect 12163 13574 12175 13626
rect 12175 13574 12189 13626
rect 12213 13574 12227 13626
rect 12227 13574 12239 13626
rect 12239 13574 12269 13626
rect 12293 13574 12303 13626
rect 12303 13574 12349 13626
rect 12053 13572 12109 13574
rect 12133 13572 12189 13574
rect 12213 13572 12269 13574
rect 12293 13572 12349 13574
rect 16492 13626 16548 13628
rect 16572 13626 16628 13628
rect 16652 13626 16708 13628
rect 16732 13626 16788 13628
rect 16492 13574 16538 13626
rect 16538 13574 16548 13626
rect 16572 13574 16602 13626
rect 16602 13574 16614 13626
rect 16614 13574 16628 13626
rect 16652 13574 16666 13626
rect 16666 13574 16678 13626
rect 16678 13574 16708 13626
rect 16732 13574 16742 13626
rect 16742 13574 16788 13626
rect 16492 13572 16548 13574
rect 16572 13572 16628 13574
rect 16652 13572 16708 13574
rect 16732 13572 16788 13574
rect 5394 13082 5450 13084
rect 5474 13082 5530 13084
rect 5554 13082 5610 13084
rect 5634 13082 5690 13084
rect 5394 13030 5440 13082
rect 5440 13030 5450 13082
rect 5474 13030 5504 13082
rect 5504 13030 5516 13082
rect 5516 13030 5530 13082
rect 5554 13030 5568 13082
rect 5568 13030 5580 13082
rect 5580 13030 5610 13082
rect 5634 13030 5644 13082
rect 5644 13030 5690 13082
rect 5394 13028 5450 13030
rect 5474 13028 5530 13030
rect 5554 13028 5610 13030
rect 5634 13028 5690 13030
rect 9833 13082 9889 13084
rect 9913 13082 9969 13084
rect 9993 13082 10049 13084
rect 10073 13082 10129 13084
rect 9833 13030 9879 13082
rect 9879 13030 9889 13082
rect 9913 13030 9943 13082
rect 9943 13030 9955 13082
rect 9955 13030 9969 13082
rect 9993 13030 10007 13082
rect 10007 13030 10019 13082
rect 10019 13030 10049 13082
rect 10073 13030 10083 13082
rect 10083 13030 10129 13082
rect 9833 13028 9889 13030
rect 9913 13028 9969 13030
rect 9993 13028 10049 13030
rect 10073 13028 10129 13030
rect 14272 13082 14328 13084
rect 14352 13082 14408 13084
rect 14432 13082 14488 13084
rect 14512 13082 14568 13084
rect 14272 13030 14318 13082
rect 14318 13030 14328 13082
rect 14352 13030 14382 13082
rect 14382 13030 14394 13082
rect 14394 13030 14408 13082
rect 14432 13030 14446 13082
rect 14446 13030 14458 13082
rect 14458 13030 14488 13082
rect 14512 13030 14522 13082
rect 14522 13030 14568 13082
rect 14272 13028 14328 13030
rect 14352 13028 14408 13030
rect 14432 13028 14488 13030
rect 14512 13028 14568 13030
rect 3175 12538 3231 12540
rect 3255 12538 3311 12540
rect 3335 12538 3391 12540
rect 3415 12538 3471 12540
rect 3175 12486 3221 12538
rect 3221 12486 3231 12538
rect 3255 12486 3285 12538
rect 3285 12486 3297 12538
rect 3297 12486 3311 12538
rect 3335 12486 3349 12538
rect 3349 12486 3361 12538
rect 3361 12486 3391 12538
rect 3415 12486 3425 12538
rect 3425 12486 3471 12538
rect 3175 12484 3231 12486
rect 3255 12484 3311 12486
rect 3335 12484 3391 12486
rect 3415 12484 3471 12486
rect 7614 12538 7670 12540
rect 7694 12538 7750 12540
rect 7774 12538 7830 12540
rect 7854 12538 7910 12540
rect 7614 12486 7660 12538
rect 7660 12486 7670 12538
rect 7694 12486 7724 12538
rect 7724 12486 7736 12538
rect 7736 12486 7750 12538
rect 7774 12486 7788 12538
rect 7788 12486 7800 12538
rect 7800 12486 7830 12538
rect 7854 12486 7864 12538
rect 7864 12486 7910 12538
rect 7614 12484 7670 12486
rect 7694 12484 7750 12486
rect 7774 12484 7830 12486
rect 7854 12484 7910 12486
rect 12053 12538 12109 12540
rect 12133 12538 12189 12540
rect 12213 12538 12269 12540
rect 12293 12538 12349 12540
rect 12053 12486 12099 12538
rect 12099 12486 12109 12538
rect 12133 12486 12163 12538
rect 12163 12486 12175 12538
rect 12175 12486 12189 12538
rect 12213 12486 12227 12538
rect 12227 12486 12239 12538
rect 12239 12486 12269 12538
rect 12293 12486 12303 12538
rect 12303 12486 12349 12538
rect 12053 12484 12109 12486
rect 12133 12484 12189 12486
rect 12213 12484 12269 12486
rect 12293 12484 12349 12486
rect 16492 12538 16548 12540
rect 16572 12538 16628 12540
rect 16652 12538 16708 12540
rect 16732 12538 16788 12540
rect 16492 12486 16538 12538
rect 16538 12486 16548 12538
rect 16572 12486 16602 12538
rect 16602 12486 16614 12538
rect 16614 12486 16628 12538
rect 16652 12486 16666 12538
rect 16666 12486 16678 12538
rect 16678 12486 16708 12538
rect 16732 12486 16742 12538
rect 16742 12486 16788 12538
rect 16492 12484 16548 12486
rect 16572 12484 16628 12486
rect 16652 12484 16708 12486
rect 16732 12484 16788 12486
rect 5394 11994 5450 11996
rect 5474 11994 5530 11996
rect 5554 11994 5610 11996
rect 5634 11994 5690 11996
rect 5394 11942 5440 11994
rect 5440 11942 5450 11994
rect 5474 11942 5504 11994
rect 5504 11942 5516 11994
rect 5516 11942 5530 11994
rect 5554 11942 5568 11994
rect 5568 11942 5580 11994
rect 5580 11942 5610 11994
rect 5634 11942 5644 11994
rect 5644 11942 5690 11994
rect 5394 11940 5450 11942
rect 5474 11940 5530 11942
rect 5554 11940 5610 11942
rect 5634 11940 5690 11942
rect 9833 11994 9889 11996
rect 9913 11994 9969 11996
rect 9993 11994 10049 11996
rect 10073 11994 10129 11996
rect 9833 11942 9879 11994
rect 9879 11942 9889 11994
rect 9913 11942 9943 11994
rect 9943 11942 9955 11994
rect 9955 11942 9969 11994
rect 9993 11942 10007 11994
rect 10007 11942 10019 11994
rect 10019 11942 10049 11994
rect 10073 11942 10083 11994
rect 10083 11942 10129 11994
rect 9833 11940 9889 11942
rect 9913 11940 9969 11942
rect 9993 11940 10049 11942
rect 10073 11940 10129 11942
rect 14272 11994 14328 11996
rect 14352 11994 14408 11996
rect 14432 11994 14488 11996
rect 14512 11994 14568 11996
rect 14272 11942 14318 11994
rect 14318 11942 14328 11994
rect 14352 11942 14382 11994
rect 14382 11942 14394 11994
rect 14394 11942 14408 11994
rect 14432 11942 14446 11994
rect 14446 11942 14458 11994
rect 14458 11942 14488 11994
rect 14512 11942 14522 11994
rect 14522 11942 14568 11994
rect 14272 11940 14328 11942
rect 14352 11940 14408 11942
rect 14432 11940 14488 11942
rect 14512 11940 14568 11942
rect 3175 11450 3231 11452
rect 3255 11450 3311 11452
rect 3335 11450 3391 11452
rect 3415 11450 3471 11452
rect 3175 11398 3221 11450
rect 3221 11398 3231 11450
rect 3255 11398 3285 11450
rect 3285 11398 3297 11450
rect 3297 11398 3311 11450
rect 3335 11398 3349 11450
rect 3349 11398 3361 11450
rect 3361 11398 3391 11450
rect 3415 11398 3425 11450
rect 3425 11398 3471 11450
rect 3175 11396 3231 11398
rect 3255 11396 3311 11398
rect 3335 11396 3391 11398
rect 3415 11396 3471 11398
rect 7614 11450 7670 11452
rect 7694 11450 7750 11452
rect 7774 11450 7830 11452
rect 7854 11450 7910 11452
rect 7614 11398 7660 11450
rect 7660 11398 7670 11450
rect 7694 11398 7724 11450
rect 7724 11398 7736 11450
rect 7736 11398 7750 11450
rect 7774 11398 7788 11450
rect 7788 11398 7800 11450
rect 7800 11398 7830 11450
rect 7854 11398 7864 11450
rect 7864 11398 7910 11450
rect 7614 11396 7670 11398
rect 7694 11396 7750 11398
rect 7774 11396 7830 11398
rect 7854 11396 7910 11398
rect 12053 11450 12109 11452
rect 12133 11450 12189 11452
rect 12213 11450 12269 11452
rect 12293 11450 12349 11452
rect 12053 11398 12099 11450
rect 12099 11398 12109 11450
rect 12133 11398 12163 11450
rect 12163 11398 12175 11450
rect 12175 11398 12189 11450
rect 12213 11398 12227 11450
rect 12227 11398 12239 11450
rect 12239 11398 12269 11450
rect 12293 11398 12303 11450
rect 12303 11398 12349 11450
rect 12053 11396 12109 11398
rect 12133 11396 12189 11398
rect 12213 11396 12269 11398
rect 12293 11396 12349 11398
rect 16492 11450 16548 11452
rect 16572 11450 16628 11452
rect 16652 11450 16708 11452
rect 16732 11450 16788 11452
rect 16492 11398 16538 11450
rect 16538 11398 16548 11450
rect 16572 11398 16602 11450
rect 16602 11398 16614 11450
rect 16614 11398 16628 11450
rect 16652 11398 16666 11450
rect 16666 11398 16678 11450
rect 16678 11398 16708 11450
rect 16732 11398 16742 11450
rect 16742 11398 16788 11450
rect 16492 11396 16548 11398
rect 16572 11396 16628 11398
rect 16652 11396 16708 11398
rect 16732 11396 16788 11398
rect 5394 10906 5450 10908
rect 5474 10906 5530 10908
rect 5554 10906 5610 10908
rect 5634 10906 5690 10908
rect 5394 10854 5440 10906
rect 5440 10854 5450 10906
rect 5474 10854 5504 10906
rect 5504 10854 5516 10906
rect 5516 10854 5530 10906
rect 5554 10854 5568 10906
rect 5568 10854 5580 10906
rect 5580 10854 5610 10906
rect 5634 10854 5644 10906
rect 5644 10854 5690 10906
rect 5394 10852 5450 10854
rect 5474 10852 5530 10854
rect 5554 10852 5610 10854
rect 5634 10852 5690 10854
rect 9833 10906 9889 10908
rect 9913 10906 9969 10908
rect 9993 10906 10049 10908
rect 10073 10906 10129 10908
rect 9833 10854 9879 10906
rect 9879 10854 9889 10906
rect 9913 10854 9943 10906
rect 9943 10854 9955 10906
rect 9955 10854 9969 10906
rect 9993 10854 10007 10906
rect 10007 10854 10019 10906
rect 10019 10854 10049 10906
rect 10073 10854 10083 10906
rect 10083 10854 10129 10906
rect 9833 10852 9889 10854
rect 9913 10852 9969 10854
rect 9993 10852 10049 10854
rect 10073 10852 10129 10854
rect 14272 10906 14328 10908
rect 14352 10906 14408 10908
rect 14432 10906 14488 10908
rect 14512 10906 14568 10908
rect 14272 10854 14318 10906
rect 14318 10854 14328 10906
rect 14352 10854 14382 10906
rect 14382 10854 14394 10906
rect 14394 10854 14408 10906
rect 14432 10854 14446 10906
rect 14446 10854 14458 10906
rect 14458 10854 14488 10906
rect 14512 10854 14522 10906
rect 14522 10854 14568 10906
rect 14272 10852 14328 10854
rect 14352 10852 14408 10854
rect 14432 10852 14488 10854
rect 14512 10852 14568 10854
rect 3175 10362 3231 10364
rect 3255 10362 3311 10364
rect 3335 10362 3391 10364
rect 3415 10362 3471 10364
rect 3175 10310 3221 10362
rect 3221 10310 3231 10362
rect 3255 10310 3285 10362
rect 3285 10310 3297 10362
rect 3297 10310 3311 10362
rect 3335 10310 3349 10362
rect 3349 10310 3361 10362
rect 3361 10310 3391 10362
rect 3415 10310 3425 10362
rect 3425 10310 3471 10362
rect 3175 10308 3231 10310
rect 3255 10308 3311 10310
rect 3335 10308 3391 10310
rect 3415 10308 3471 10310
rect 7614 10362 7670 10364
rect 7694 10362 7750 10364
rect 7774 10362 7830 10364
rect 7854 10362 7910 10364
rect 7614 10310 7660 10362
rect 7660 10310 7670 10362
rect 7694 10310 7724 10362
rect 7724 10310 7736 10362
rect 7736 10310 7750 10362
rect 7774 10310 7788 10362
rect 7788 10310 7800 10362
rect 7800 10310 7830 10362
rect 7854 10310 7864 10362
rect 7864 10310 7910 10362
rect 7614 10308 7670 10310
rect 7694 10308 7750 10310
rect 7774 10308 7830 10310
rect 7854 10308 7910 10310
rect 12053 10362 12109 10364
rect 12133 10362 12189 10364
rect 12213 10362 12269 10364
rect 12293 10362 12349 10364
rect 12053 10310 12099 10362
rect 12099 10310 12109 10362
rect 12133 10310 12163 10362
rect 12163 10310 12175 10362
rect 12175 10310 12189 10362
rect 12213 10310 12227 10362
rect 12227 10310 12239 10362
rect 12239 10310 12269 10362
rect 12293 10310 12303 10362
rect 12303 10310 12349 10362
rect 12053 10308 12109 10310
rect 12133 10308 12189 10310
rect 12213 10308 12269 10310
rect 12293 10308 12349 10310
rect 16492 10362 16548 10364
rect 16572 10362 16628 10364
rect 16652 10362 16708 10364
rect 16732 10362 16788 10364
rect 16492 10310 16538 10362
rect 16538 10310 16548 10362
rect 16572 10310 16602 10362
rect 16602 10310 16614 10362
rect 16614 10310 16628 10362
rect 16652 10310 16666 10362
rect 16666 10310 16678 10362
rect 16678 10310 16708 10362
rect 16732 10310 16742 10362
rect 16742 10310 16788 10362
rect 16492 10308 16548 10310
rect 16572 10308 16628 10310
rect 16652 10308 16708 10310
rect 16732 10308 16788 10310
rect 5394 9818 5450 9820
rect 5474 9818 5530 9820
rect 5554 9818 5610 9820
rect 5634 9818 5690 9820
rect 5394 9766 5440 9818
rect 5440 9766 5450 9818
rect 5474 9766 5504 9818
rect 5504 9766 5516 9818
rect 5516 9766 5530 9818
rect 5554 9766 5568 9818
rect 5568 9766 5580 9818
rect 5580 9766 5610 9818
rect 5634 9766 5644 9818
rect 5644 9766 5690 9818
rect 5394 9764 5450 9766
rect 5474 9764 5530 9766
rect 5554 9764 5610 9766
rect 5634 9764 5690 9766
rect 9833 9818 9889 9820
rect 9913 9818 9969 9820
rect 9993 9818 10049 9820
rect 10073 9818 10129 9820
rect 9833 9766 9879 9818
rect 9879 9766 9889 9818
rect 9913 9766 9943 9818
rect 9943 9766 9955 9818
rect 9955 9766 9969 9818
rect 9993 9766 10007 9818
rect 10007 9766 10019 9818
rect 10019 9766 10049 9818
rect 10073 9766 10083 9818
rect 10083 9766 10129 9818
rect 9833 9764 9889 9766
rect 9913 9764 9969 9766
rect 9993 9764 10049 9766
rect 10073 9764 10129 9766
rect 14272 9818 14328 9820
rect 14352 9818 14408 9820
rect 14432 9818 14488 9820
rect 14512 9818 14568 9820
rect 14272 9766 14318 9818
rect 14318 9766 14328 9818
rect 14352 9766 14382 9818
rect 14382 9766 14394 9818
rect 14394 9766 14408 9818
rect 14432 9766 14446 9818
rect 14446 9766 14458 9818
rect 14458 9766 14488 9818
rect 14512 9766 14522 9818
rect 14522 9766 14568 9818
rect 14272 9764 14328 9766
rect 14352 9764 14408 9766
rect 14432 9764 14488 9766
rect 14512 9764 14568 9766
rect 3175 9274 3231 9276
rect 3255 9274 3311 9276
rect 3335 9274 3391 9276
rect 3415 9274 3471 9276
rect 3175 9222 3221 9274
rect 3221 9222 3231 9274
rect 3255 9222 3285 9274
rect 3285 9222 3297 9274
rect 3297 9222 3311 9274
rect 3335 9222 3349 9274
rect 3349 9222 3361 9274
rect 3361 9222 3391 9274
rect 3415 9222 3425 9274
rect 3425 9222 3471 9274
rect 3175 9220 3231 9222
rect 3255 9220 3311 9222
rect 3335 9220 3391 9222
rect 3415 9220 3471 9222
rect 7614 9274 7670 9276
rect 7694 9274 7750 9276
rect 7774 9274 7830 9276
rect 7854 9274 7910 9276
rect 7614 9222 7660 9274
rect 7660 9222 7670 9274
rect 7694 9222 7724 9274
rect 7724 9222 7736 9274
rect 7736 9222 7750 9274
rect 7774 9222 7788 9274
rect 7788 9222 7800 9274
rect 7800 9222 7830 9274
rect 7854 9222 7864 9274
rect 7864 9222 7910 9274
rect 7614 9220 7670 9222
rect 7694 9220 7750 9222
rect 7774 9220 7830 9222
rect 7854 9220 7910 9222
rect 12053 9274 12109 9276
rect 12133 9274 12189 9276
rect 12213 9274 12269 9276
rect 12293 9274 12349 9276
rect 12053 9222 12099 9274
rect 12099 9222 12109 9274
rect 12133 9222 12163 9274
rect 12163 9222 12175 9274
rect 12175 9222 12189 9274
rect 12213 9222 12227 9274
rect 12227 9222 12239 9274
rect 12239 9222 12269 9274
rect 12293 9222 12303 9274
rect 12303 9222 12349 9274
rect 12053 9220 12109 9222
rect 12133 9220 12189 9222
rect 12213 9220 12269 9222
rect 12293 9220 12349 9222
rect 16492 9274 16548 9276
rect 16572 9274 16628 9276
rect 16652 9274 16708 9276
rect 16732 9274 16788 9276
rect 16492 9222 16538 9274
rect 16538 9222 16548 9274
rect 16572 9222 16602 9274
rect 16602 9222 16614 9274
rect 16614 9222 16628 9274
rect 16652 9222 16666 9274
rect 16666 9222 16678 9274
rect 16678 9222 16708 9274
rect 16732 9222 16742 9274
rect 16742 9222 16788 9274
rect 16492 9220 16548 9222
rect 16572 9220 16628 9222
rect 16652 9220 16708 9222
rect 16732 9220 16788 9222
rect 5394 8730 5450 8732
rect 5474 8730 5530 8732
rect 5554 8730 5610 8732
rect 5634 8730 5690 8732
rect 5394 8678 5440 8730
rect 5440 8678 5450 8730
rect 5474 8678 5504 8730
rect 5504 8678 5516 8730
rect 5516 8678 5530 8730
rect 5554 8678 5568 8730
rect 5568 8678 5580 8730
rect 5580 8678 5610 8730
rect 5634 8678 5644 8730
rect 5644 8678 5690 8730
rect 5394 8676 5450 8678
rect 5474 8676 5530 8678
rect 5554 8676 5610 8678
rect 5634 8676 5690 8678
rect 9833 8730 9889 8732
rect 9913 8730 9969 8732
rect 9993 8730 10049 8732
rect 10073 8730 10129 8732
rect 9833 8678 9879 8730
rect 9879 8678 9889 8730
rect 9913 8678 9943 8730
rect 9943 8678 9955 8730
rect 9955 8678 9969 8730
rect 9993 8678 10007 8730
rect 10007 8678 10019 8730
rect 10019 8678 10049 8730
rect 10073 8678 10083 8730
rect 10083 8678 10129 8730
rect 9833 8676 9889 8678
rect 9913 8676 9969 8678
rect 9993 8676 10049 8678
rect 10073 8676 10129 8678
rect 14272 8730 14328 8732
rect 14352 8730 14408 8732
rect 14432 8730 14488 8732
rect 14512 8730 14568 8732
rect 14272 8678 14318 8730
rect 14318 8678 14328 8730
rect 14352 8678 14382 8730
rect 14382 8678 14394 8730
rect 14394 8678 14408 8730
rect 14432 8678 14446 8730
rect 14446 8678 14458 8730
rect 14458 8678 14488 8730
rect 14512 8678 14522 8730
rect 14522 8678 14568 8730
rect 14272 8676 14328 8678
rect 14352 8676 14408 8678
rect 14432 8676 14488 8678
rect 14512 8676 14568 8678
rect 3175 8186 3231 8188
rect 3255 8186 3311 8188
rect 3335 8186 3391 8188
rect 3415 8186 3471 8188
rect 3175 8134 3221 8186
rect 3221 8134 3231 8186
rect 3255 8134 3285 8186
rect 3285 8134 3297 8186
rect 3297 8134 3311 8186
rect 3335 8134 3349 8186
rect 3349 8134 3361 8186
rect 3361 8134 3391 8186
rect 3415 8134 3425 8186
rect 3425 8134 3471 8186
rect 3175 8132 3231 8134
rect 3255 8132 3311 8134
rect 3335 8132 3391 8134
rect 3415 8132 3471 8134
rect 7614 8186 7670 8188
rect 7694 8186 7750 8188
rect 7774 8186 7830 8188
rect 7854 8186 7910 8188
rect 7614 8134 7660 8186
rect 7660 8134 7670 8186
rect 7694 8134 7724 8186
rect 7724 8134 7736 8186
rect 7736 8134 7750 8186
rect 7774 8134 7788 8186
rect 7788 8134 7800 8186
rect 7800 8134 7830 8186
rect 7854 8134 7864 8186
rect 7864 8134 7910 8186
rect 7614 8132 7670 8134
rect 7694 8132 7750 8134
rect 7774 8132 7830 8134
rect 7854 8132 7910 8134
rect 12053 8186 12109 8188
rect 12133 8186 12189 8188
rect 12213 8186 12269 8188
rect 12293 8186 12349 8188
rect 12053 8134 12099 8186
rect 12099 8134 12109 8186
rect 12133 8134 12163 8186
rect 12163 8134 12175 8186
rect 12175 8134 12189 8186
rect 12213 8134 12227 8186
rect 12227 8134 12239 8186
rect 12239 8134 12269 8186
rect 12293 8134 12303 8186
rect 12303 8134 12349 8186
rect 12053 8132 12109 8134
rect 12133 8132 12189 8134
rect 12213 8132 12269 8134
rect 12293 8132 12349 8134
rect 5394 7642 5450 7644
rect 5474 7642 5530 7644
rect 5554 7642 5610 7644
rect 5634 7642 5690 7644
rect 5394 7590 5440 7642
rect 5440 7590 5450 7642
rect 5474 7590 5504 7642
rect 5504 7590 5516 7642
rect 5516 7590 5530 7642
rect 5554 7590 5568 7642
rect 5568 7590 5580 7642
rect 5580 7590 5610 7642
rect 5634 7590 5644 7642
rect 5644 7590 5690 7642
rect 5394 7588 5450 7590
rect 5474 7588 5530 7590
rect 5554 7588 5610 7590
rect 5634 7588 5690 7590
rect 9833 7642 9889 7644
rect 9913 7642 9969 7644
rect 9993 7642 10049 7644
rect 10073 7642 10129 7644
rect 9833 7590 9879 7642
rect 9879 7590 9889 7642
rect 9913 7590 9943 7642
rect 9943 7590 9955 7642
rect 9955 7590 9969 7642
rect 9993 7590 10007 7642
rect 10007 7590 10019 7642
rect 10019 7590 10049 7642
rect 10073 7590 10083 7642
rect 10083 7590 10129 7642
rect 9833 7588 9889 7590
rect 9913 7588 9969 7590
rect 9993 7588 10049 7590
rect 10073 7588 10129 7590
rect 14272 7642 14328 7644
rect 14352 7642 14408 7644
rect 14432 7642 14488 7644
rect 14512 7642 14568 7644
rect 14272 7590 14318 7642
rect 14318 7590 14328 7642
rect 14352 7590 14382 7642
rect 14382 7590 14394 7642
rect 14394 7590 14408 7642
rect 14432 7590 14446 7642
rect 14446 7590 14458 7642
rect 14458 7590 14488 7642
rect 14512 7590 14522 7642
rect 14522 7590 14568 7642
rect 14272 7588 14328 7590
rect 14352 7588 14408 7590
rect 14432 7588 14488 7590
rect 14512 7588 14568 7590
rect 3175 7098 3231 7100
rect 3255 7098 3311 7100
rect 3335 7098 3391 7100
rect 3415 7098 3471 7100
rect 3175 7046 3221 7098
rect 3221 7046 3231 7098
rect 3255 7046 3285 7098
rect 3285 7046 3297 7098
rect 3297 7046 3311 7098
rect 3335 7046 3349 7098
rect 3349 7046 3361 7098
rect 3361 7046 3391 7098
rect 3415 7046 3425 7098
rect 3425 7046 3471 7098
rect 3175 7044 3231 7046
rect 3255 7044 3311 7046
rect 3335 7044 3391 7046
rect 3415 7044 3471 7046
rect 7614 7098 7670 7100
rect 7694 7098 7750 7100
rect 7774 7098 7830 7100
rect 7854 7098 7910 7100
rect 7614 7046 7660 7098
rect 7660 7046 7670 7098
rect 7694 7046 7724 7098
rect 7724 7046 7736 7098
rect 7736 7046 7750 7098
rect 7774 7046 7788 7098
rect 7788 7046 7800 7098
rect 7800 7046 7830 7098
rect 7854 7046 7864 7098
rect 7864 7046 7910 7098
rect 7614 7044 7670 7046
rect 7694 7044 7750 7046
rect 7774 7044 7830 7046
rect 7854 7044 7910 7046
rect 12053 7098 12109 7100
rect 12133 7098 12189 7100
rect 12213 7098 12269 7100
rect 12293 7098 12349 7100
rect 12053 7046 12099 7098
rect 12099 7046 12109 7098
rect 12133 7046 12163 7098
rect 12163 7046 12175 7098
rect 12175 7046 12189 7098
rect 12213 7046 12227 7098
rect 12227 7046 12239 7098
rect 12239 7046 12269 7098
rect 12293 7046 12303 7098
rect 12303 7046 12349 7098
rect 12053 7044 12109 7046
rect 12133 7044 12189 7046
rect 12213 7044 12269 7046
rect 12293 7044 12349 7046
rect 16492 8186 16548 8188
rect 16572 8186 16628 8188
rect 16652 8186 16708 8188
rect 16732 8186 16788 8188
rect 16492 8134 16538 8186
rect 16538 8134 16548 8186
rect 16572 8134 16602 8186
rect 16602 8134 16614 8186
rect 16614 8134 16628 8186
rect 16652 8134 16666 8186
rect 16666 8134 16678 8186
rect 16678 8134 16708 8186
rect 16732 8134 16742 8186
rect 16742 8134 16788 8186
rect 16492 8132 16548 8134
rect 16572 8132 16628 8134
rect 16652 8132 16708 8134
rect 16732 8132 16788 8134
rect 5394 6554 5450 6556
rect 5474 6554 5530 6556
rect 5554 6554 5610 6556
rect 5634 6554 5690 6556
rect 5394 6502 5440 6554
rect 5440 6502 5450 6554
rect 5474 6502 5504 6554
rect 5504 6502 5516 6554
rect 5516 6502 5530 6554
rect 5554 6502 5568 6554
rect 5568 6502 5580 6554
rect 5580 6502 5610 6554
rect 5634 6502 5644 6554
rect 5644 6502 5690 6554
rect 5394 6500 5450 6502
rect 5474 6500 5530 6502
rect 5554 6500 5610 6502
rect 5634 6500 5690 6502
rect 9833 6554 9889 6556
rect 9913 6554 9969 6556
rect 9993 6554 10049 6556
rect 10073 6554 10129 6556
rect 9833 6502 9879 6554
rect 9879 6502 9889 6554
rect 9913 6502 9943 6554
rect 9943 6502 9955 6554
rect 9955 6502 9969 6554
rect 9993 6502 10007 6554
rect 10007 6502 10019 6554
rect 10019 6502 10049 6554
rect 10073 6502 10083 6554
rect 10083 6502 10129 6554
rect 9833 6500 9889 6502
rect 9913 6500 9969 6502
rect 9993 6500 10049 6502
rect 10073 6500 10129 6502
rect 14272 6554 14328 6556
rect 14352 6554 14408 6556
rect 14432 6554 14488 6556
rect 14512 6554 14568 6556
rect 14272 6502 14318 6554
rect 14318 6502 14328 6554
rect 14352 6502 14382 6554
rect 14382 6502 14394 6554
rect 14394 6502 14408 6554
rect 14432 6502 14446 6554
rect 14446 6502 14458 6554
rect 14458 6502 14488 6554
rect 14512 6502 14522 6554
rect 14522 6502 14568 6554
rect 14272 6500 14328 6502
rect 14352 6500 14408 6502
rect 14432 6500 14488 6502
rect 14512 6500 14568 6502
rect 3175 6010 3231 6012
rect 3255 6010 3311 6012
rect 3335 6010 3391 6012
rect 3415 6010 3471 6012
rect 3175 5958 3221 6010
rect 3221 5958 3231 6010
rect 3255 5958 3285 6010
rect 3285 5958 3297 6010
rect 3297 5958 3311 6010
rect 3335 5958 3349 6010
rect 3349 5958 3361 6010
rect 3361 5958 3391 6010
rect 3415 5958 3425 6010
rect 3425 5958 3471 6010
rect 3175 5956 3231 5958
rect 3255 5956 3311 5958
rect 3335 5956 3391 5958
rect 3415 5956 3471 5958
rect 7614 6010 7670 6012
rect 7694 6010 7750 6012
rect 7774 6010 7830 6012
rect 7854 6010 7910 6012
rect 7614 5958 7660 6010
rect 7660 5958 7670 6010
rect 7694 5958 7724 6010
rect 7724 5958 7736 6010
rect 7736 5958 7750 6010
rect 7774 5958 7788 6010
rect 7788 5958 7800 6010
rect 7800 5958 7830 6010
rect 7854 5958 7864 6010
rect 7864 5958 7910 6010
rect 7614 5956 7670 5958
rect 7694 5956 7750 5958
rect 7774 5956 7830 5958
rect 7854 5956 7910 5958
rect 12053 6010 12109 6012
rect 12133 6010 12189 6012
rect 12213 6010 12269 6012
rect 12293 6010 12349 6012
rect 12053 5958 12099 6010
rect 12099 5958 12109 6010
rect 12133 5958 12163 6010
rect 12163 5958 12175 6010
rect 12175 5958 12189 6010
rect 12213 5958 12227 6010
rect 12227 5958 12239 6010
rect 12239 5958 12269 6010
rect 12293 5958 12303 6010
rect 12303 5958 12349 6010
rect 12053 5956 12109 5958
rect 12133 5956 12189 5958
rect 12213 5956 12269 5958
rect 12293 5956 12349 5958
rect 5394 5466 5450 5468
rect 5474 5466 5530 5468
rect 5554 5466 5610 5468
rect 5634 5466 5690 5468
rect 5394 5414 5440 5466
rect 5440 5414 5450 5466
rect 5474 5414 5504 5466
rect 5504 5414 5516 5466
rect 5516 5414 5530 5466
rect 5554 5414 5568 5466
rect 5568 5414 5580 5466
rect 5580 5414 5610 5466
rect 5634 5414 5644 5466
rect 5644 5414 5690 5466
rect 5394 5412 5450 5414
rect 5474 5412 5530 5414
rect 5554 5412 5610 5414
rect 5634 5412 5690 5414
rect 9833 5466 9889 5468
rect 9913 5466 9969 5468
rect 9993 5466 10049 5468
rect 10073 5466 10129 5468
rect 9833 5414 9879 5466
rect 9879 5414 9889 5466
rect 9913 5414 9943 5466
rect 9943 5414 9955 5466
rect 9955 5414 9969 5466
rect 9993 5414 10007 5466
rect 10007 5414 10019 5466
rect 10019 5414 10049 5466
rect 10073 5414 10083 5466
rect 10083 5414 10129 5466
rect 9833 5412 9889 5414
rect 9913 5412 9969 5414
rect 9993 5412 10049 5414
rect 10073 5412 10129 5414
rect 14272 5466 14328 5468
rect 14352 5466 14408 5468
rect 14432 5466 14488 5468
rect 14512 5466 14568 5468
rect 14272 5414 14318 5466
rect 14318 5414 14328 5466
rect 14352 5414 14382 5466
rect 14382 5414 14394 5466
rect 14394 5414 14408 5466
rect 14432 5414 14446 5466
rect 14446 5414 14458 5466
rect 14458 5414 14488 5466
rect 14512 5414 14522 5466
rect 14522 5414 14568 5466
rect 14272 5412 14328 5414
rect 14352 5412 14408 5414
rect 14432 5412 14488 5414
rect 14512 5412 14568 5414
rect 18711 40282 18767 40284
rect 18791 40282 18847 40284
rect 18871 40282 18927 40284
rect 18951 40282 19007 40284
rect 18711 40230 18757 40282
rect 18757 40230 18767 40282
rect 18791 40230 18821 40282
rect 18821 40230 18833 40282
rect 18833 40230 18847 40282
rect 18871 40230 18885 40282
rect 18885 40230 18897 40282
rect 18897 40230 18927 40282
rect 18951 40230 18961 40282
rect 18961 40230 19007 40282
rect 18711 40228 18767 40230
rect 18791 40228 18847 40230
rect 18871 40228 18927 40230
rect 18951 40228 19007 40230
rect 18711 39194 18767 39196
rect 18791 39194 18847 39196
rect 18871 39194 18927 39196
rect 18951 39194 19007 39196
rect 18711 39142 18757 39194
rect 18757 39142 18767 39194
rect 18791 39142 18821 39194
rect 18821 39142 18833 39194
rect 18833 39142 18847 39194
rect 18871 39142 18885 39194
rect 18885 39142 18897 39194
rect 18897 39142 18927 39194
rect 18951 39142 18961 39194
rect 18961 39142 19007 39194
rect 18711 39140 18767 39142
rect 18791 39140 18847 39142
rect 18871 39140 18927 39142
rect 18951 39140 19007 39142
rect 18711 38106 18767 38108
rect 18791 38106 18847 38108
rect 18871 38106 18927 38108
rect 18951 38106 19007 38108
rect 18711 38054 18757 38106
rect 18757 38054 18767 38106
rect 18791 38054 18821 38106
rect 18821 38054 18833 38106
rect 18833 38054 18847 38106
rect 18871 38054 18885 38106
rect 18885 38054 18897 38106
rect 18897 38054 18927 38106
rect 18951 38054 18961 38106
rect 18961 38054 19007 38106
rect 18711 38052 18767 38054
rect 18791 38052 18847 38054
rect 18871 38052 18927 38054
rect 18951 38052 19007 38054
rect 18711 37018 18767 37020
rect 18791 37018 18847 37020
rect 18871 37018 18927 37020
rect 18951 37018 19007 37020
rect 18711 36966 18757 37018
rect 18757 36966 18767 37018
rect 18791 36966 18821 37018
rect 18821 36966 18833 37018
rect 18833 36966 18847 37018
rect 18871 36966 18885 37018
rect 18885 36966 18897 37018
rect 18897 36966 18927 37018
rect 18951 36966 18961 37018
rect 18961 36966 19007 37018
rect 18711 36964 18767 36966
rect 18791 36964 18847 36966
rect 18871 36964 18927 36966
rect 18951 36964 19007 36966
rect 18711 35930 18767 35932
rect 18791 35930 18847 35932
rect 18871 35930 18927 35932
rect 18951 35930 19007 35932
rect 18711 35878 18757 35930
rect 18757 35878 18767 35930
rect 18791 35878 18821 35930
rect 18821 35878 18833 35930
rect 18833 35878 18847 35930
rect 18871 35878 18885 35930
rect 18885 35878 18897 35930
rect 18897 35878 18927 35930
rect 18951 35878 18961 35930
rect 18961 35878 19007 35930
rect 18711 35876 18767 35878
rect 18791 35876 18847 35878
rect 18871 35876 18927 35878
rect 18951 35876 19007 35878
rect 18711 34842 18767 34844
rect 18791 34842 18847 34844
rect 18871 34842 18927 34844
rect 18951 34842 19007 34844
rect 18711 34790 18757 34842
rect 18757 34790 18767 34842
rect 18791 34790 18821 34842
rect 18821 34790 18833 34842
rect 18833 34790 18847 34842
rect 18871 34790 18885 34842
rect 18885 34790 18897 34842
rect 18897 34790 18927 34842
rect 18951 34790 18961 34842
rect 18961 34790 19007 34842
rect 18711 34788 18767 34790
rect 18791 34788 18847 34790
rect 18871 34788 18927 34790
rect 18951 34788 19007 34790
rect 18510 34348 18512 34368
rect 18512 34348 18564 34368
rect 18564 34348 18566 34368
rect 18510 34312 18566 34348
rect 18711 33754 18767 33756
rect 18791 33754 18847 33756
rect 18871 33754 18927 33756
rect 18951 33754 19007 33756
rect 18711 33702 18757 33754
rect 18757 33702 18767 33754
rect 18791 33702 18821 33754
rect 18821 33702 18833 33754
rect 18833 33702 18847 33754
rect 18871 33702 18885 33754
rect 18885 33702 18897 33754
rect 18897 33702 18927 33754
rect 18951 33702 18961 33754
rect 18961 33702 19007 33754
rect 18711 33700 18767 33702
rect 18791 33700 18847 33702
rect 18871 33700 18927 33702
rect 18951 33700 19007 33702
rect 18711 32666 18767 32668
rect 18791 32666 18847 32668
rect 18871 32666 18927 32668
rect 18951 32666 19007 32668
rect 18711 32614 18757 32666
rect 18757 32614 18767 32666
rect 18791 32614 18821 32666
rect 18821 32614 18833 32666
rect 18833 32614 18847 32666
rect 18871 32614 18885 32666
rect 18885 32614 18897 32666
rect 18897 32614 18927 32666
rect 18951 32614 18961 32666
rect 18961 32614 19007 32666
rect 18711 32612 18767 32614
rect 18791 32612 18847 32614
rect 18871 32612 18927 32614
rect 18951 32612 19007 32614
rect 18711 31578 18767 31580
rect 18791 31578 18847 31580
rect 18871 31578 18927 31580
rect 18951 31578 19007 31580
rect 18711 31526 18757 31578
rect 18757 31526 18767 31578
rect 18791 31526 18821 31578
rect 18821 31526 18833 31578
rect 18833 31526 18847 31578
rect 18871 31526 18885 31578
rect 18885 31526 18897 31578
rect 18897 31526 18927 31578
rect 18951 31526 18961 31578
rect 18961 31526 19007 31578
rect 18711 31524 18767 31526
rect 18791 31524 18847 31526
rect 18871 31524 18927 31526
rect 18951 31524 19007 31526
rect 18711 30490 18767 30492
rect 18791 30490 18847 30492
rect 18871 30490 18927 30492
rect 18951 30490 19007 30492
rect 18711 30438 18757 30490
rect 18757 30438 18767 30490
rect 18791 30438 18821 30490
rect 18821 30438 18833 30490
rect 18833 30438 18847 30490
rect 18871 30438 18885 30490
rect 18885 30438 18897 30490
rect 18897 30438 18927 30490
rect 18951 30438 18961 30490
rect 18961 30438 19007 30490
rect 18711 30436 18767 30438
rect 18791 30436 18847 30438
rect 18871 30436 18927 30438
rect 18951 30436 19007 30438
rect 18711 29402 18767 29404
rect 18791 29402 18847 29404
rect 18871 29402 18927 29404
rect 18951 29402 19007 29404
rect 18711 29350 18757 29402
rect 18757 29350 18767 29402
rect 18791 29350 18821 29402
rect 18821 29350 18833 29402
rect 18833 29350 18847 29402
rect 18871 29350 18885 29402
rect 18885 29350 18897 29402
rect 18897 29350 18927 29402
rect 18951 29350 18961 29402
rect 18961 29350 19007 29402
rect 18711 29348 18767 29350
rect 18791 29348 18847 29350
rect 18871 29348 18927 29350
rect 18951 29348 19007 29350
rect 18711 28314 18767 28316
rect 18791 28314 18847 28316
rect 18871 28314 18927 28316
rect 18951 28314 19007 28316
rect 18711 28262 18757 28314
rect 18757 28262 18767 28314
rect 18791 28262 18821 28314
rect 18821 28262 18833 28314
rect 18833 28262 18847 28314
rect 18871 28262 18885 28314
rect 18885 28262 18897 28314
rect 18897 28262 18927 28314
rect 18951 28262 18961 28314
rect 18961 28262 19007 28314
rect 18711 28260 18767 28262
rect 18791 28260 18847 28262
rect 18871 28260 18927 28262
rect 18951 28260 19007 28262
rect 18602 28056 18658 28112
rect 18711 27226 18767 27228
rect 18791 27226 18847 27228
rect 18871 27226 18927 27228
rect 18951 27226 19007 27228
rect 18711 27174 18757 27226
rect 18757 27174 18767 27226
rect 18791 27174 18821 27226
rect 18821 27174 18833 27226
rect 18833 27174 18847 27226
rect 18871 27174 18885 27226
rect 18885 27174 18897 27226
rect 18897 27174 18927 27226
rect 18951 27174 18961 27226
rect 18961 27174 19007 27226
rect 18711 27172 18767 27174
rect 18791 27172 18847 27174
rect 18871 27172 18927 27174
rect 18951 27172 19007 27174
rect 18711 26138 18767 26140
rect 18791 26138 18847 26140
rect 18871 26138 18927 26140
rect 18951 26138 19007 26140
rect 18711 26086 18757 26138
rect 18757 26086 18767 26138
rect 18791 26086 18821 26138
rect 18821 26086 18833 26138
rect 18833 26086 18847 26138
rect 18871 26086 18885 26138
rect 18885 26086 18897 26138
rect 18897 26086 18927 26138
rect 18951 26086 18961 26138
rect 18961 26086 19007 26138
rect 18711 26084 18767 26086
rect 18791 26084 18847 26086
rect 18871 26084 18927 26086
rect 18951 26084 19007 26086
rect 18711 25050 18767 25052
rect 18791 25050 18847 25052
rect 18871 25050 18927 25052
rect 18951 25050 19007 25052
rect 18711 24998 18757 25050
rect 18757 24998 18767 25050
rect 18791 24998 18821 25050
rect 18821 24998 18833 25050
rect 18833 24998 18847 25050
rect 18871 24998 18885 25050
rect 18885 24998 18897 25050
rect 18897 24998 18927 25050
rect 18951 24998 18961 25050
rect 18961 24998 19007 25050
rect 18711 24996 18767 24998
rect 18791 24996 18847 24998
rect 18871 24996 18927 24998
rect 18951 24996 19007 24998
rect 18326 15544 18382 15600
rect 18711 23962 18767 23964
rect 18791 23962 18847 23964
rect 18871 23962 18927 23964
rect 18951 23962 19007 23964
rect 18711 23910 18757 23962
rect 18757 23910 18767 23962
rect 18791 23910 18821 23962
rect 18821 23910 18833 23962
rect 18833 23910 18847 23962
rect 18871 23910 18885 23962
rect 18885 23910 18897 23962
rect 18897 23910 18927 23962
rect 18951 23910 18961 23962
rect 18961 23910 19007 23962
rect 18711 23908 18767 23910
rect 18791 23908 18847 23910
rect 18871 23908 18927 23910
rect 18951 23908 19007 23910
rect 18711 22874 18767 22876
rect 18791 22874 18847 22876
rect 18871 22874 18927 22876
rect 18951 22874 19007 22876
rect 18711 22822 18757 22874
rect 18757 22822 18767 22874
rect 18791 22822 18821 22874
rect 18821 22822 18833 22874
rect 18833 22822 18847 22874
rect 18871 22822 18885 22874
rect 18885 22822 18897 22874
rect 18897 22822 18927 22874
rect 18951 22822 18961 22874
rect 18961 22822 19007 22874
rect 18711 22820 18767 22822
rect 18791 22820 18847 22822
rect 18871 22820 18927 22822
rect 18951 22820 19007 22822
rect 18510 22072 18566 22128
rect 18711 21786 18767 21788
rect 18791 21786 18847 21788
rect 18871 21786 18927 21788
rect 18951 21786 19007 21788
rect 18711 21734 18757 21786
rect 18757 21734 18767 21786
rect 18791 21734 18821 21786
rect 18821 21734 18833 21786
rect 18833 21734 18847 21786
rect 18871 21734 18885 21786
rect 18885 21734 18897 21786
rect 18897 21734 18927 21786
rect 18951 21734 18961 21786
rect 18961 21734 19007 21786
rect 18711 21732 18767 21734
rect 18791 21732 18847 21734
rect 18871 21732 18927 21734
rect 18951 21732 19007 21734
rect 18711 20698 18767 20700
rect 18791 20698 18847 20700
rect 18871 20698 18927 20700
rect 18951 20698 19007 20700
rect 18711 20646 18757 20698
rect 18757 20646 18767 20698
rect 18791 20646 18821 20698
rect 18821 20646 18833 20698
rect 18833 20646 18847 20698
rect 18871 20646 18885 20698
rect 18885 20646 18897 20698
rect 18897 20646 18927 20698
rect 18951 20646 18961 20698
rect 18961 20646 19007 20698
rect 18711 20644 18767 20646
rect 18791 20644 18847 20646
rect 18871 20644 18927 20646
rect 18951 20644 19007 20646
rect 18711 19610 18767 19612
rect 18791 19610 18847 19612
rect 18871 19610 18927 19612
rect 18951 19610 19007 19612
rect 18711 19558 18757 19610
rect 18757 19558 18767 19610
rect 18791 19558 18821 19610
rect 18821 19558 18833 19610
rect 18833 19558 18847 19610
rect 18871 19558 18885 19610
rect 18885 19558 18897 19610
rect 18897 19558 18927 19610
rect 18951 19558 18961 19610
rect 18961 19558 19007 19610
rect 18711 19556 18767 19558
rect 18791 19556 18847 19558
rect 18871 19556 18927 19558
rect 18951 19556 19007 19558
rect 18711 18522 18767 18524
rect 18791 18522 18847 18524
rect 18871 18522 18927 18524
rect 18951 18522 19007 18524
rect 18711 18470 18757 18522
rect 18757 18470 18767 18522
rect 18791 18470 18821 18522
rect 18821 18470 18833 18522
rect 18833 18470 18847 18522
rect 18871 18470 18885 18522
rect 18885 18470 18897 18522
rect 18897 18470 18927 18522
rect 18951 18470 18961 18522
rect 18961 18470 19007 18522
rect 18711 18468 18767 18470
rect 18791 18468 18847 18470
rect 18871 18468 18927 18470
rect 18951 18468 19007 18470
rect 18711 17434 18767 17436
rect 18791 17434 18847 17436
rect 18871 17434 18927 17436
rect 18951 17434 19007 17436
rect 18711 17382 18757 17434
rect 18757 17382 18767 17434
rect 18791 17382 18821 17434
rect 18821 17382 18833 17434
rect 18833 17382 18847 17434
rect 18871 17382 18885 17434
rect 18885 17382 18897 17434
rect 18897 17382 18927 17434
rect 18951 17382 18961 17434
rect 18961 17382 19007 17434
rect 18711 17380 18767 17382
rect 18791 17380 18847 17382
rect 18871 17380 18927 17382
rect 18951 17380 19007 17382
rect 18711 16346 18767 16348
rect 18791 16346 18847 16348
rect 18871 16346 18927 16348
rect 18951 16346 19007 16348
rect 18711 16294 18757 16346
rect 18757 16294 18767 16346
rect 18791 16294 18821 16346
rect 18821 16294 18833 16346
rect 18833 16294 18847 16346
rect 18871 16294 18885 16346
rect 18885 16294 18897 16346
rect 18897 16294 18927 16346
rect 18951 16294 18961 16346
rect 18961 16294 19007 16346
rect 18711 16292 18767 16294
rect 18791 16292 18847 16294
rect 18871 16292 18927 16294
rect 18951 16292 19007 16294
rect 18711 15258 18767 15260
rect 18791 15258 18847 15260
rect 18871 15258 18927 15260
rect 18951 15258 19007 15260
rect 18711 15206 18757 15258
rect 18757 15206 18767 15258
rect 18791 15206 18821 15258
rect 18821 15206 18833 15258
rect 18833 15206 18847 15258
rect 18871 15206 18885 15258
rect 18885 15206 18897 15258
rect 18897 15206 18927 15258
rect 18951 15206 18961 15258
rect 18961 15206 19007 15258
rect 18711 15204 18767 15206
rect 18791 15204 18847 15206
rect 18871 15204 18927 15206
rect 18951 15204 19007 15206
rect 18711 14170 18767 14172
rect 18791 14170 18847 14172
rect 18871 14170 18927 14172
rect 18951 14170 19007 14172
rect 18711 14118 18757 14170
rect 18757 14118 18767 14170
rect 18791 14118 18821 14170
rect 18821 14118 18833 14170
rect 18833 14118 18847 14170
rect 18871 14118 18885 14170
rect 18885 14118 18897 14170
rect 18897 14118 18927 14170
rect 18951 14118 18961 14170
rect 18961 14118 19007 14170
rect 18711 14116 18767 14118
rect 18791 14116 18847 14118
rect 18871 14116 18927 14118
rect 18951 14116 19007 14118
rect 18711 13082 18767 13084
rect 18791 13082 18847 13084
rect 18871 13082 18927 13084
rect 18951 13082 19007 13084
rect 18711 13030 18757 13082
rect 18757 13030 18767 13082
rect 18791 13030 18821 13082
rect 18821 13030 18833 13082
rect 18833 13030 18847 13082
rect 18871 13030 18885 13082
rect 18885 13030 18897 13082
rect 18897 13030 18927 13082
rect 18951 13030 18961 13082
rect 18961 13030 19007 13082
rect 18711 13028 18767 13030
rect 18791 13028 18847 13030
rect 18871 13028 18927 13030
rect 18951 13028 19007 13030
rect 18711 11994 18767 11996
rect 18791 11994 18847 11996
rect 18871 11994 18927 11996
rect 18951 11994 19007 11996
rect 18711 11942 18757 11994
rect 18757 11942 18767 11994
rect 18791 11942 18821 11994
rect 18821 11942 18833 11994
rect 18833 11942 18847 11994
rect 18871 11942 18885 11994
rect 18885 11942 18897 11994
rect 18897 11942 18927 11994
rect 18951 11942 18961 11994
rect 18961 11942 19007 11994
rect 18711 11940 18767 11942
rect 18791 11940 18847 11942
rect 18871 11940 18927 11942
rect 18951 11940 19007 11942
rect 18711 10906 18767 10908
rect 18791 10906 18847 10908
rect 18871 10906 18927 10908
rect 18951 10906 19007 10908
rect 18711 10854 18757 10906
rect 18757 10854 18767 10906
rect 18791 10854 18821 10906
rect 18821 10854 18833 10906
rect 18833 10854 18847 10906
rect 18871 10854 18885 10906
rect 18885 10854 18897 10906
rect 18897 10854 18927 10906
rect 18951 10854 18961 10906
rect 18961 10854 19007 10906
rect 18711 10852 18767 10854
rect 18791 10852 18847 10854
rect 18871 10852 18927 10854
rect 18951 10852 19007 10854
rect 18711 9818 18767 9820
rect 18791 9818 18847 9820
rect 18871 9818 18927 9820
rect 18951 9818 19007 9820
rect 18711 9766 18757 9818
rect 18757 9766 18767 9818
rect 18791 9766 18821 9818
rect 18821 9766 18833 9818
rect 18833 9766 18847 9818
rect 18871 9766 18885 9818
rect 18885 9766 18897 9818
rect 18897 9766 18927 9818
rect 18951 9766 18961 9818
rect 18961 9766 19007 9818
rect 18711 9764 18767 9766
rect 18791 9764 18847 9766
rect 18871 9764 18927 9766
rect 18951 9764 19007 9766
rect 18510 9324 18512 9344
rect 18512 9324 18564 9344
rect 18564 9324 18566 9344
rect 18510 9288 18566 9324
rect 18711 8730 18767 8732
rect 18791 8730 18847 8732
rect 18871 8730 18927 8732
rect 18951 8730 19007 8732
rect 18711 8678 18757 8730
rect 18757 8678 18767 8730
rect 18791 8678 18821 8730
rect 18821 8678 18833 8730
rect 18833 8678 18847 8730
rect 18871 8678 18885 8730
rect 18885 8678 18897 8730
rect 18897 8678 18927 8730
rect 18951 8678 18961 8730
rect 18961 8678 19007 8730
rect 18711 8676 18767 8678
rect 18791 8676 18847 8678
rect 18871 8676 18927 8678
rect 18951 8676 19007 8678
rect 16492 7098 16548 7100
rect 16572 7098 16628 7100
rect 16652 7098 16708 7100
rect 16732 7098 16788 7100
rect 16492 7046 16538 7098
rect 16538 7046 16548 7098
rect 16572 7046 16602 7098
rect 16602 7046 16614 7098
rect 16614 7046 16628 7098
rect 16652 7046 16666 7098
rect 16666 7046 16678 7098
rect 16678 7046 16708 7098
rect 16732 7046 16742 7098
rect 16742 7046 16788 7098
rect 16492 7044 16548 7046
rect 16572 7044 16628 7046
rect 16652 7044 16708 7046
rect 16732 7044 16788 7046
rect 16492 6010 16548 6012
rect 16572 6010 16628 6012
rect 16652 6010 16708 6012
rect 16732 6010 16788 6012
rect 16492 5958 16538 6010
rect 16538 5958 16548 6010
rect 16572 5958 16602 6010
rect 16602 5958 16614 6010
rect 16614 5958 16628 6010
rect 16652 5958 16666 6010
rect 16666 5958 16678 6010
rect 16678 5958 16708 6010
rect 16732 5958 16742 6010
rect 16742 5958 16788 6010
rect 16492 5956 16548 5958
rect 16572 5956 16628 5958
rect 16652 5956 16708 5958
rect 16732 5956 16788 5958
rect 3175 4922 3231 4924
rect 3255 4922 3311 4924
rect 3335 4922 3391 4924
rect 3415 4922 3471 4924
rect 3175 4870 3221 4922
rect 3221 4870 3231 4922
rect 3255 4870 3285 4922
rect 3285 4870 3297 4922
rect 3297 4870 3311 4922
rect 3335 4870 3349 4922
rect 3349 4870 3361 4922
rect 3361 4870 3391 4922
rect 3415 4870 3425 4922
rect 3425 4870 3471 4922
rect 3175 4868 3231 4870
rect 3255 4868 3311 4870
rect 3335 4868 3391 4870
rect 3415 4868 3471 4870
rect 7614 4922 7670 4924
rect 7694 4922 7750 4924
rect 7774 4922 7830 4924
rect 7854 4922 7910 4924
rect 7614 4870 7660 4922
rect 7660 4870 7670 4922
rect 7694 4870 7724 4922
rect 7724 4870 7736 4922
rect 7736 4870 7750 4922
rect 7774 4870 7788 4922
rect 7788 4870 7800 4922
rect 7800 4870 7830 4922
rect 7854 4870 7864 4922
rect 7864 4870 7910 4922
rect 7614 4868 7670 4870
rect 7694 4868 7750 4870
rect 7774 4868 7830 4870
rect 7854 4868 7910 4870
rect 12053 4922 12109 4924
rect 12133 4922 12189 4924
rect 12213 4922 12269 4924
rect 12293 4922 12349 4924
rect 12053 4870 12099 4922
rect 12099 4870 12109 4922
rect 12133 4870 12163 4922
rect 12163 4870 12175 4922
rect 12175 4870 12189 4922
rect 12213 4870 12227 4922
rect 12227 4870 12239 4922
rect 12239 4870 12269 4922
rect 12293 4870 12303 4922
rect 12303 4870 12349 4922
rect 12053 4868 12109 4870
rect 12133 4868 12189 4870
rect 12213 4868 12269 4870
rect 12293 4868 12349 4870
rect 5394 4378 5450 4380
rect 5474 4378 5530 4380
rect 5554 4378 5610 4380
rect 5634 4378 5690 4380
rect 5394 4326 5440 4378
rect 5440 4326 5450 4378
rect 5474 4326 5504 4378
rect 5504 4326 5516 4378
rect 5516 4326 5530 4378
rect 5554 4326 5568 4378
rect 5568 4326 5580 4378
rect 5580 4326 5610 4378
rect 5634 4326 5644 4378
rect 5644 4326 5690 4378
rect 5394 4324 5450 4326
rect 5474 4324 5530 4326
rect 5554 4324 5610 4326
rect 5634 4324 5690 4326
rect 9833 4378 9889 4380
rect 9913 4378 9969 4380
rect 9993 4378 10049 4380
rect 10073 4378 10129 4380
rect 9833 4326 9879 4378
rect 9879 4326 9889 4378
rect 9913 4326 9943 4378
rect 9943 4326 9955 4378
rect 9955 4326 9969 4378
rect 9993 4326 10007 4378
rect 10007 4326 10019 4378
rect 10019 4326 10049 4378
rect 10073 4326 10083 4378
rect 10083 4326 10129 4378
rect 9833 4324 9889 4326
rect 9913 4324 9969 4326
rect 9993 4324 10049 4326
rect 10073 4324 10129 4326
rect 14272 4378 14328 4380
rect 14352 4378 14408 4380
rect 14432 4378 14488 4380
rect 14512 4378 14568 4380
rect 14272 4326 14318 4378
rect 14318 4326 14328 4378
rect 14352 4326 14382 4378
rect 14382 4326 14394 4378
rect 14394 4326 14408 4378
rect 14432 4326 14446 4378
rect 14446 4326 14458 4378
rect 14458 4326 14488 4378
rect 14512 4326 14522 4378
rect 14522 4326 14568 4378
rect 14272 4324 14328 4326
rect 14352 4324 14408 4326
rect 14432 4324 14488 4326
rect 14512 4324 14568 4326
rect 3175 3834 3231 3836
rect 3255 3834 3311 3836
rect 3335 3834 3391 3836
rect 3415 3834 3471 3836
rect 3175 3782 3221 3834
rect 3221 3782 3231 3834
rect 3255 3782 3285 3834
rect 3285 3782 3297 3834
rect 3297 3782 3311 3834
rect 3335 3782 3349 3834
rect 3349 3782 3361 3834
rect 3361 3782 3391 3834
rect 3415 3782 3425 3834
rect 3425 3782 3471 3834
rect 3175 3780 3231 3782
rect 3255 3780 3311 3782
rect 3335 3780 3391 3782
rect 3415 3780 3471 3782
rect 7614 3834 7670 3836
rect 7694 3834 7750 3836
rect 7774 3834 7830 3836
rect 7854 3834 7910 3836
rect 7614 3782 7660 3834
rect 7660 3782 7670 3834
rect 7694 3782 7724 3834
rect 7724 3782 7736 3834
rect 7736 3782 7750 3834
rect 7774 3782 7788 3834
rect 7788 3782 7800 3834
rect 7800 3782 7830 3834
rect 7854 3782 7864 3834
rect 7864 3782 7910 3834
rect 7614 3780 7670 3782
rect 7694 3780 7750 3782
rect 7774 3780 7830 3782
rect 7854 3780 7910 3782
rect 12053 3834 12109 3836
rect 12133 3834 12189 3836
rect 12213 3834 12269 3836
rect 12293 3834 12349 3836
rect 12053 3782 12099 3834
rect 12099 3782 12109 3834
rect 12133 3782 12163 3834
rect 12163 3782 12175 3834
rect 12175 3782 12189 3834
rect 12213 3782 12227 3834
rect 12227 3782 12239 3834
rect 12239 3782 12269 3834
rect 12293 3782 12303 3834
rect 12303 3782 12349 3834
rect 12053 3780 12109 3782
rect 12133 3780 12189 3782
rect 12213 3780 12269 3782
rect 12293 3780 12349 3782
rect 3175 2746 3231 2748
rect 3255 2746 3311 2748
rect 3335 2746 3391 2748
rect 3415 2746 3471 2748
rect 3175 2694 3221 2746
rect 3221 2694 3231 2746
rect 3255 2694 3285 2746
rect 3285 2694 3297 2746
rect 3297 2694 3311 2746
rect 3335 2694 3349 2746
rect 3349 2694 3361 2746
rect 3361 2694 3391 2746
rect 3415 2694 3425 2746
rect 3425 2694 3471 2746
rect 3175 2692 3231 2694
rect 3255 2692 3311 2694
rect 3335 2692 3391 2694
rect 3415 2692 3471 2694
rect 5394 3290 5450 3292
rect 5474 3290 5530 3292
rect 5554 3290 5610 3292
rect 5634 3290 5690 3292
rect 5394 3238 5440 3290
rect 5440 3238 5450 3290
rect 5474 3238 5504 3290
rect 5504 3238 5516 3290
rect 5516 3238 5530 3290
rect 5554 3238 5568 3290
rect 5568 3238 5580 3290
rect 5580 3238 5610 3290
rect 5634 3238 5644 3290
rect 5644 3238 5690 3290
rect 5394 3236 5450 3238
rect 5474 3236 5530 3238
rect 5554 3236 5610 3238
rect 5634 3236 5690 3238
rect 9833 3290 9889 3292
rect 9913 3290 9969 3292
rect 9993 3290 10049 3292
rect 10073 3290 10129 3292
rect 9833 3238 9879 3290
rect 9879 3238 9889 3290
rect 9913 3238 9943 3290
rect 9943 3238 9955 3290
rect 9955 3238 9969 3290
rect 9993 3238 10007 3290
rect 10007 3238 10019 3290
rect 10019 3238 10049 3290
rect 10073 3238 10083 3290
rect 10083 3238 10129 3290
rect 9833 3236 9889 3238
rect 9913 3236 9969 3238
rect 9993 3236 10049 3238
rect 10073 3236 10129 3238
rect 14272 3290 14328 3292
rect 14352 3290 14408 3292
rect 14432 3290 14488 3292
rect 14512 3290 14568 3292
rect 14272 3238 14318 3290
rect 14318 3238 14328 3290
rect 14352 3238 14382 3290
rect 14382 3238 14394 3290
rect 14394 3238 14408 3290
rect 14432 3238 14446 3290
rect 14446 3238 14458 3290
rect 14458 3238 14488 3290
rect 14512 3238 14522 3290
rect 14522 3238 14568 3290
rect 14272 3236 14328 3238
rect 14352 3236 14408 3238
rect 14432 3236 14488 3238
rect 14512 3236 14568 3238
rect 16492 4922 16548 4924
rect 16572 4922 16628 4924
rect 16652 4922 16708 4924
rect 16732 4922 16788 4924
rect 16492 4870 16538 4922
rect 16538 4870 16548 4922
rect 16572 4870 16602 4922
rect 16602 4870 16614 4922
rect 16614 4870 16628 4922
rect 16652 4870 16666 4922
rect 16666 4870 16678 4922
rect 16678 4870 16708 4922
rect 16732 4870 16742 4922
rect 16742 4870 16788 4922
rect 16492 4868 16548 4870
rect 16572 4868 16628 4870
rect 16652 4868 16708 4870
rect 16732 4868 16788 4870
rect 16492 3834 16548 3836
rect 16572 3834 16628 3836
rect 16652 3834 16708 3836
rect 16732 3834 16788 3836
rect 16492 3782 16538 3834
rect 16538 3782 16548 3834
rect 16572 3782 16602 3834
rect 16602 3782 16614 3834
rect 16614 3782 16628 3834
rect 16652 3782 16666 3834
rect 16666 3782 16678 3834
rect 16678 3782 16708 3834
rect 16732 3782 16742 3834
rect 16742 3782 16788 3834
rect 16492 3780 16548 3782
rect 16572 3780 16628 3782
rect 16652 3780 16708 3782
rect 16732 3780 16788 3782
rect 18711 7642 18767 7644
rect 18791 7642 18847 7644
rect 18871 7642 18927 7644
rect 18951 7642 19007 7644
rect 18711 7590 18757 7642
rect 18757 7590 18767 7642
rect 18791 7590 18821 7642
rect 18821 7590 18833 7642
rect 18833 7590 18847 7642
rect 18871 7590 18885 7642
rect 18885 7590 18897 7642
rect 18897 7590 18927 7642
rect 18951 7590 18961 7642
rect 18961 7590 19007 7642
rect 18711 7588 18767 7590
rect 18791 7588 18847 7590
rect 18871 7588 18927 7590
rect 18951 7588 19007 7590
rect 18711 6554 18767 6556
rect 18791 6554 18847 6556
rect 18871 6554 18927 6556
rect 18951 6554 19007 6556
rect 18711 6502 18757 6554
rect 18757 6502 18767 6554
rect 18791 6502 18821 6554
rect 18821 6502 18833 6554
rect 18833 6502 18847 6554
rect 18871 6502 18885 6554
rect 18885 6502 18897 6554
rect 18897 6502 18927 6554
rect 18951 6502 18961 6554
rect 18961 6502 19007 6554
rect 18711 6500 18767 6502
rect 18791 6500 18847 6502
rect 18871 6500 18927 6502
rect 18951 6500 19007 6502
rect 18711 5466 18767 5468
rect 18791 5466 18847 5468
rect 18871 5466 18927 5468
rect 18951 5466 19007 5468
rect 18711 5414 18757 5466
rect 18757 5414 18767 5466
rect 18791 5414 18821 5466
rect 18821 5414 18833 5466
rect 18833 5414 18847 5466
rect 18871 5414 18885 5466
rect 18885 5414 18897 5466
rect 18897 5414 18927 5466
rect 18951 5414 18961 5466
rect 18961 5414 19007 5466
rect 18711 5412 18767 5414
rect 18791 5412 18847 5414
rect 18871 5412 18927 5414
rect 18951 5412 19007 5414
rect 18711 4378 18767 4380
rect 18791 4378 18847 4380
rect 18871 4378 18927 4380
rect 18951 4378 19007 4380
rect 18711 4326 18757 4378
rect 18757 4326 18767 4378
rect 18791 4326 18821 4378
rect 18821 4326 18833 4378
rect 18833 4326 18847 4378
rect 18871 4326 18885 4378
rect 18885 4326 18897 4378
rect 18897 4326 18927 4378
rect 18951 4326 18961 4378
rect 18961 4326 19007 4378
rect 18711 4324 18767 4326
rect 18791 4324 18847 4326
rect 18871 4324 18927 4326
rect 18951 4324 19007 4326
rect 7614 2746 7670 2748
rect 7694 2746 7750 2748
rect 7774 2746 7830 2748
rect 7854 2746 7910 2748
rect 7614 2694 7660 2746
rect 7660 2694 7670 2746
rect 7694 2694 7724 2746
rect 7724 2694 7736 2746
rect 7736 2694 7750 2746
rect 7774 2694 7788 2746
rect 7788 2694 7800 2746
rect 7800 2694 7830 2746
rect 7854 2694 7864 2746
rect 7864 2694 7910 2746
rect 7614 2692 7670 2694
rect 7694 2692 7750 2694
rect 7774 2692 7830 2694
rect 7854 2692 7910 2694
rect 12053 2746 12109 2748
rect 12133 2746 12189 2748
rect 12213 2746 12269 2748
rect 12293 2746 12349 2748
rect 12053 2694 12099 2746
rect 12099 2694 12109 2746
rect 12133 2694 12163 2746
rect 12163 2694 12175 2746
rect 12175 2694 12189 2746
rect 12213 2694 12227 2746
rect 12227 2694 12239 2746
rect 12239 2694 12269 2746
rect 12293 2694 12303 2746
rect 12303 2694 12349 2746
rect 12053 2692 12109 2694
rect 12133 2692 12189 2694
rect 12213 2692 12269 2694
rect 12293 2692 12349 2694
rect 16492 2746 16548 2748
rect 16572 2746 16628 2748
rect 16652 2746 16708 2748
rect 16732 2746 16788 2748
rect 16492 2694 16538 2746
rect 16538 2694 16548 2746
rect 16572 2694 16602 2746
rect 16602 2694 16614 2746
rect 16614 2694 16628 2746
rect 16652 2694 16666 2746
rect 16666 2694 16678 2746
rect 16678 2694 16708 2746
rect 16732 2694 16742 2746
rect 16742 2694 16788 2746
rect 16492 2692 16548 2694
rect 16572 2692 16628 2694
rect 16652 2692 16708 2694
rect 16732 2692 16788 2694
rect 18326 3032 18382 3088
rect 18711 3290 18767 3292
rect 18791 3290 18847 3292
rect 18871 3290 18927 3292
rect 18951 3290 19007 3292
rect 18711 3238 18757 3290
rect 18757 3238 18767 3290
rect 18791 3238 18821 3290
rect 18821 3238 18833 3290
rect 18833 3238 18847 3290
rect 18871 3238 18885 3290
rect 18885 3238 18897 3290
rect 18897 3238 18927 3290
rect 18951 3238 18961 3290
rect 18961 3238 19007 3290
rect 18711 3236 18767 3238
rect 18791 3236 18847 3238
rect 18871 3236 18927 3238
rect 18951 3236 19007 3238
rect 5394 2202 5450 2204
rect 5474 2202 5530 2204
rect 5554 2202 5610 2204
rect 5634 2202 5690 2204
rect 5394 2150 5440 2202
rect 5440 2150 5450 2202
rect 5474 2150 5504 2202
rect 5504 2150 5516 2202
rect 5516 2150 5530 2202
rect 5554 2150 5568 2202
rect 5568 2150 5580 2202
rect 5580 2150 5610 2202
rect 5634 2150 5644 2202
rect 5644 2150 5690 2202
rect 5394 2148 5450 2150
rect 5474 2148 5530 2150
rect 5554 2148 5610 2150
rect 5634 2148 5690 2150
rect 9833 2202 9889 2204
rect 9913 2202 9969 2204
rect 9993 2202 10049 2204
rect 10073 2202 10129 2204
rect 9833 2150 9879 2202
rect 9879 2150 9889 2202
rect 9913 2150 9943 2202
rect 9943 2150 9955 2202
rect 9955 2150 9969 2202
rect 9993 2150 10007 2202
rect 10007 2150 10019 2202
rect 10019 2150 10049 2202
rect 10073 2150 10083 2202
rect 10083 2150 10129 2202
rect 9833 2148 9889 2150
rect 9913 2148 9969 2150
rect 9993 2148 10049 2150
rect 10073 2148 10129 2150
rect 14272 2202 14328 2204
rect 14352 2202 14408 2204
rect 14432 2202 14488 2204
rect 14512 2202 14568 2204
rect 14272 2150 14318 2202
rect 14318 2150 14328 2202
rect 14352 2150 14382 2202
rect 14382 2150 14394 2202
rect 14394 2150 14408 2202
rect 14432 2150 14446 2202
rect 14446 2150 14458 2202
rect 14458 2150 14488 2202
rect 14512 2150 14522 2202
rect 14522 2150 14568 2202
rect 14272 2148 14328 2150
rect 14352 2148 14408 2150
rect 14432 2148 14488 2150
rect 14512 2148 14568 2150
rect 18711 2202 18767 2204
rect 18791 2202 18847 2204
rect 18871 2202 18927 2204
rect 18951 2202 19007 2204
rect 18711 2150 18757 2202
rect 18757 2150 18767 2202
rect 18791 2150 18821 2202
rect 18821 2150 18833 2202
rect 18833 2150 18847 2202
rect 18871 2150 18885 2202
rect 18885 2150 18897 2202
rect 18897 2150 18927 2202
rect 18951 2150 18961 2202
rect 18961 2150 19007 2202
rect 18711 2148 18767 2150
rect 18791 2148 18847 2150
rect 18871 2148 18927 2150
rect 18951 2148 19007 2150
<< metal3 >>
rect 3165 47360 3481 47361
rect 3165 47296 3171 47360
rect 3235 47296 3251 47360
rect 3315 47296 3331 47360
rect 3395 47296 3411 47360
rect 3475 47296 3481 47360
rect 3165 47295 3481 47296
rect 7604 47360 7920 47361
rect 7604 47296 7610 47360
rect 7674 47296 7690 47360
rect 7754 47296 7770 47360
rect 7834 47296 7850 47360
rect 7914 47296 7920 47360
rect 7604 47295 7920 47296
rect 12043 47360 12359 47361
rect 12043 47296 12049 47360
rect 12113 47296 12129 47360
rect 12193 47296 12209 47360
rect 12273 47296 12289 47360
rect 12353 47296 12359 47360
rect 12043 47295 12359 47296
rect 16482 47360 16798 47361
rect 16482 47296 16488 47360
rect 16552 47296 16568 47360
rect 16632 47296 16648 47360
rect 16712 47296 16728 47360
rect 16792 47296 16798 47360
rect 16482 47295 16798 47296
rect 18505 47154 18571 47157
rect 18505 47152 19626 47154
rect 18505 47096 18510 47152
rect 18566 47096 19626 47152
rect 18505 47094 19626 47096
rect 18505 47091 18571 47094
rect 19566 46912 19626 47094
rect 5384 46816 5700 46817
rect 5384 46752 5390 46816
rect 5454 46752 5470 46816
rect 5534 46752 5550 46816
rect 5614 46752 5630 46816
rect 5694 46752 5700 46816
rect 5384 46751 5700 46752
rect 9823 46816 10139 46817
rect 9823 46752 9829 46816
rect 9893 46752 9909 46816
rect 9973 46752 9989 46816
rect 10053 46752 10069 46816
rect 10133 46752 10139 46816
rect 9823 46751 10139 46752
rect 14262 46816 14578 46817
rect 14262 46752 14268 46816
rect 14332 46752 14348 46816
rect 14412 46752 14428 46816
rect 14492 46752 14508 46816
rect 14572 46752 14578 46816
rect 14262 46751 14578 46752
rect 18701 46816 19017 46817
rect 18701 46752 18707 46816
rect 18771 46752 18787 46816
rect 18851 46752 18867 46816
rect 18931 46752 18947 46816
rect 19011 46752 19017 46816
rect 19200 46792 20000 46912
rect 18701 46751 19017 46752
rect 3165 46272 3481 46273
rect 3165 46208 3171 46272
rect 3235 46208 3251 46272
rect 3315 46208 3331 46272
rect 3395 46208 3411 46272
rect 3475 46208 3481 46272
rect 3165 46207 3481 46208
rect 7604 46272 7920 46273
rect 7604 46208 7610 46272
rect 7674 46208 7690 46272
rect 7754 46208 7770 46272
rect 7834 46208 7850 46272
rect 7914 46208 7920 46272
rect 7604 46207 7920 46208
rect 12043 46272 12359 46273
rect 12043 46208 12049 46272
rect 12113 46208 12129 46272
rect 12193 46208 12209 46272
rect 12273 46208 12289 46272
rect 12353 46208 12359 46272
rect 12043 46207 12359 46208
rect 16482 46272 16798 46273
rect 16482 46208 16488 46272
rect 16552 46208 16568 46272
rect 16632 46208 16648 46272
rect 16712 46208 16728 46272
rect 16792 46208 16798 46272
rect 16482 46207 16798 46208
rect 5384 45728 5700 45729
rect 5384 45664 5390 45728
rect 5454 45664 5470 45728
rect 5534 45664 5550 45728
rect 5614 45664 5630 45728
rect 5694 45664 5700 45728
rect 5384 45663 5700 45664
rect 9823 45728 10139 45729
rect 9823 45664 9829 45728
rect 9893 45664 9909 45728
rect 9973 45664 9989 45728
rect 10053 45664 10069 45728
rect 10133 45664 10139 45728
rect 9823 45663 10139 45664
rect 14262 45728 14578 45729
rect 14262 45664 14268 45728
rect 14332 45664 14348 45728
rect 14412 45664 14428 45728
rect 14492 45664 14508 45728
rect 14572 45664 14578 45728
rect 14262 45663 14578 45664
rect 18701 45728 19017 45729
rect 18701 45664 18707 45728
rect 18771 45664 18787 45728
rect 18851 45664 18867 45728
rect 18931 45664 18947 45728
rect 19011 45664 19017 45728
rect 18701 45663 19017 45664
rect 3165 45184 3481 45185
rect 3165 45120 3171 45184
rect 3235 45120 3251 45184
rect 3315 45120 3331 45184
rect 3395 45120 3411 45184
rect 3475 45120 3481 45184
rect 3165 45119 3481 45120
rect 7604 45184 7920 45185
rect 7604 45120 7610 45184
rect 7674 45120 7690 45184
rect 7754 45120 7770 45184
rect 7834 45120 7850 45184
rect 7914 45120 7920 45184
rect 7604 45119 7920 45120
rect 12043 45184 12359 45185
rect 12043 45120 12049 45184
rect 12113 45120 12129 45184
rect 12193 45120 12209 45184
rect 12273 45120 12289 45184
rect 12353 45120 12359 45184
rect 12043 45119 12359 45120
rect 16482 45184 16798 45185
rect 16482 45120 16488 45184
rect 16552 45120 16568 45184
rect 16632 45120 16648 45184
rect 16712 45120 16728 45184
rect 16792 45120 16798 45184
rect 16482 45119 16798 45120
rect 5384 44640 5700 44641
rect 5384 44576 5390 44640
rect 5454 44576 5470 44640
rect 5534 44576 5550 44640
rect 5614 44576 5630 44640
rect 5694 44576 5700 44640
rect 5384 44575 5700 44576
rect 9823 44640 10139 44641
rect 9823 44576 9829 44640
rect 9893 44576 9909 44640
rect 9973 44576 9989 44640
rect 10053 44576 10069 44640
rect 10133 44576 10139 44640
rect 9823 44575 10139 44576
rect 14262 44640 14578 44641
rect 14262 44576 14268 44640
rect 14332 44576 14348 44640
rect 14412 44576 14428 44640
rect 14492 44576 14508 44640
rect 14572 44576 14578 44640
rect 14262 44575 14578 44576
rect 18701 44640 19017 44641
rect 18701 44576 18707 44640
rect 18771 44576 18787 44640
rect 18851 44576 18867 44640
rect 18931 44576 18947 44640
rect 19011 44576 19017 44640
rect 18701 44575 19017 44576
rect 3165 44096 3481 44097
rect 3165 44032 3171 44096
rect 3235 44032 3251 44096
rect 3315 44032 3331 44096
rect 3395 44032 3411 44096
rect 3475 44032 3481 44096
rect 3165 44031 3481 44032
rect 7604 44096 7920 44097
rect 7604 44032 7610 44096
rect 7674 44032 7690 44096
rect 7754 44032 7770 44096
rect 7834 44032 7850 44096
rect 7914 44032 7920 44096
rect 7604 44031 7920 44032
rect 12043 44096 12359 44097
rect 12043 44032 12049 44096
rect 12113 44032 12129 44096
rect 12193 44032 12209 44096
rect 12273 44032 12289 44096
rect 12353 44032 12359 44096
rect 12043 44031 12359 44032
rect 16482 44096 16798 44097
rect 16482 44032 16488 44096
rect 16552 44032 16568 44096
rect 16632 44032 16648 44096
rect 16712 44032 16728 44096
rect 16792 44032 16798 44096
rect 16482 44031 16798 44032
rect 5384 43552 5700 43553
rect 5384 43488 5390 43552
rect 5454 43488 5470 43552
rect 5534 43488 5550 43552
rect 5614 43488 5630 43552
rect 5694 43488 5700 43552
rect 5384 43487 5700 43488
rect 9823 43552 10139 43553
rect 9823 43488 9829 43552
rect 9893 43488 9909 43552
rect 9973 43488 9989 43552
rect 10053 43488 10069 43552
rect 10133 43488 10139 43552
rect 9823 43487 10139 43488
rect 14262 43552 14578 43553
rect 14262 43488 14268 43552
rect 14332 43488 14348 43552
rect 14412 43488 14428 43552
rect 14492 43488 14508 43552
rect 14572 43488 14578 43552
rect 14262 43487 14578 43488
rect 18701 43552 19017 43553
rect 18701 43488 18707 43552
rect 18771 43488 18787 43552
rect 18851 43488 18867 43552
rect 18931 43488 18947 43552
rect 19011 43488 19017 43552
rect 18701 43487 19017 43488
rect 3165 43008 3481 43009
rect 3165 42944 3171 43008
rect 3235 42944 3251 43008
rect 3315 42944 3331 43008
rect 3395 42944 3411 43008
rect 3475 42944 3481 43008
rect 3165 42943 3481 42944
rect 7604 43008 7920 43009
rect 7604 42944 7610 43008
rect 7674 42944 7690 43008
rect 7754 42944 7770 43008
rect 7834 42944 7850 43008
rect 7914 42944 7920 43008
rect 7604 42943 7920 42944
rect 12043 43008 12359 43009
rect 12043 42944 12049 43008
rect 12113 42944 12129 43008
rect 12193 42944 12209 43008
rect 12273 42944 12289 43008
rect 12353 42944 12359 43008
rect 12043 42943 12359 42944
rect 16482 43008 16798 43009
rect 16482 42944 16488 43008
rect 16552 42944 16568 43008
rect 16632 42944 16648 43008
rect 16712 42944 16728 43008
rect 16792 42944 16798 43008
rect 16482 42943 16798 42944
rect 5384 42464 5700 42465
rect 5384 42400 5390 42464
rect 5454 42400 5470 42464
rect 5534 42400 5550 42464
rect 5614 42400 5630 42464
rect 5694 42400 5700 42464
rect 5384 42399 5700 42400
rect 9823 42464 10139 42465
rect 9823 42400 9829 42464
rect 9893 42400 9909 42464
rect 9973 42400 9989 42464
rect 10053 42400 10069 42464
rect 10133 42400 10139 42464
rect 9823 42399 10139 42400
rect 14262 42464 14578 42465
rect 14262 42400 14268 42464
rect 14332 42400 14348 42464
rect 14412 42400 14428 42464
rect 14492 42400 14508 42464
rect 14572 42400 14578 42464
rect 14262 42399 14578 42400
rect 18701 42464 19017 42465
rect 18701 42400 18707 42464
rect 18771 42400 18787 42464
rect 18851 42400 18867 42464
rect 18931 42400 18947 42464
rect 19011 42400 19017 42464
rect 18701 42399 19017 42400
rect 3165 41920 3481 41921
rect 3165 41856 3171 41920
rect 3235 41856 3251 41920
rect 3315 41856 3331 41920
rect 3395 41856 3411 41920
rect 3475 41856 3481 41920
rect 3165 41855 3481 41856
rect 7604 41920 7920 41921
rect 7604 41856 7610 41920
rect 7674 41856 7690 41920
rect 7754 41856 7770 41920
rect 7834 41856 7850 41920
rect 7914 41856 7920 41920
rect 7604 41855 7920 41856
rect 12043 41920 12359 41921
rect 12043 41856 12049 41920
rect 12113 41856 12129 41920
rect 12193 41856 12209 41920
rect 12273 41856 12289 41920
rect 12353 41856 12359 41920
rect 12043 41855 12359 41856
rect 16482 41920 16798 41921
rect 16482 41856 16488 41920
rect 16552 41856 16568 41920
rect 16632 41856 16648 41920
rect 16712 41856 16728 41920
rect 16792 41856 16798 41920
rect 16482 41855 16798 41856
rect 5384 41376 5700 41377
rect 5384 41312 5390 41376
rect 5454 41312 5470 41376
rect 5534 41312 5550 41376
rect 5614 41312 5630 41376
rect 5694 41312 5700 41376
rect 5384 41311 5700 41312
rect 9823 41376 10139 41377
rect 9823 41312 9829 41376
rect 9893 41312 9909 41376
rect 9973 41312 9989 41376
rect 10053 41312 10069 41376
rect 10133 41312 10139 41376
rect 9823 41311 10139 41312
rect 14262 41376 14578 41377
rect 14262 41312 14268 41376
rect 14332 41312 14348 41376
rect 14412 41312 14428 41376
rect 14492 41312 14508 41376
rect 14572 41312 14578 41376
rect 14262 41311 14578 41312
rect 18701 41376 19017 41377
rect 18701 41312 18707 41376
rect 18771 41312 18787 41376
rect 18851 41312 18867 41376
rect 18931 41312 18947 41376
rect 19011 41312 19017 41376
rect 18701 41311 19017 41312
rect 3165 40832 3481 40833
rect 3165 40768 3171 40832
rect 3235 40768 3251 40832
rect 3315 40768 3331 40832
rect 3395 40768 3411 40832
rect 3475 40768 3481 40832
rect 3165 40767 3481 40768
rect 7604 40832 7920 40833
rect 7604 40768 7610 40832
rect 7674 40768 7690 40832
rect 7754 40768 7770 40832
rect 7834 40768 7850 40832
rect 7914 40768 7920 40832
rect 7604 40767 7920 40768
rect 12043 40832 12359 40833
rect 12043 40768 12049 40832
rect 12113 40768 12129 40832
rect 12193 40768 12209 40832
rect 12273 40768 12289 40832
rect 12353 40768 12359 40832
rect 12043 40767 12359 40768
rect 16482 40832 16798 40833
rect 16482 40768 16488 40832
rect 16552 40768 16568 40832
rect 16632 40768 16648 40832
rect 16712 40768 16728 40832
rect 16792 40768 16798 40832
rect 16482 40767 16798 40768
rect 18045 40626 18111 40629
rect 19200 40626 20000 40656
rect 18045 40624 20000 40626
rect 18045 40568 18050 40624
rect 18106 40568 20000 40624
rect 18045 40566 20000 40568
rect 18045 40563 18111 40566
rect 19200 40536 20000 40566
rect 5384 40288 5700 40289
rect 5384 40224 5390 40288
rect 5454 40224 5470 40288
rect 5534 40224 5550 40288
rect 5614 40224 5630 40288
rect 5694 40224 5700 40288
rect 5384 40223 5700 40224
rect 9823 40288 10139 40289
rect 9823 40224 9829 40288
rect 9893 40224 9909 40288
rect 9973 40224 9989 40288
rect 10053 40224 10069 40288
rect 10133 40224 10139 40288
rect 9823 40223 10139 40224
rect 14262 40288 14578 40289
rect 14262 40224 14268 40288
rect 14332 40224 14348 40288
rect 14412 40224 14428 40288
rect 14492 40224 14508 40288
rect 14572 40224 14578 40288
rect 14262 40223 14578 40224
rect 18701 40288 19017 40289
rect 18701 40224 18707 40288
rect 18771 40224 18787 40288
rect 18851 40224 18867 40288
rect 18931 40224 18947 40288
rect 19011 40224 19017 40288
rect 18701 40223 19017 40224
rect 3165 39744 3481 39745
rect 3165 39680 3171 39744
rect 3235 39680 3251 39744
rect 3315 39680 3331 39744
rect 3395 39680 3411 39744
rect 3475 39680 3481 39744
rect 3165 39679 3481 39680
rect 7604 39744 7920 39745
rect 7604 39680 7610 39744
rect 7674 39680 7690 39744
rect 7754 39680 7770 39744
rect 7834 39680 7850 39744
rect 7914 39680 7920 39744
rect 7604 39679 7920 39680
rect 12043 39744 12359 39745
rect 12043 39680 12049 39744
rect 12113 39680 12129 39744
rect 12193 39680 12209 39744
rect 12273 39680 12289 39744
rect 12353 39680 12359 39744
rect 12043 39679 12359 39680
rect 16482 39744 16798 39745
rect 16482 39680 16488 39744
rect 16552 39680 16568 39744
rect 16632 39680 16648 39744
rect 16712 39680 16728 39744
rect 16792 39680 16798 39744
rect 16482 39679 16798 39680
rect 5384 39200 5700 39201
rect 5384 39136 5390 39200
rect 5454 39136 5470 39200
rect 5534 39136 5550 39200
rect 5614 39136 5630 39200
rect 5694 39136 5700 39200
rect 5384 39135 5700 39136
rect 9823 39200 10139 39201
rect 9823 39136 9829 39200
rect 9893 39136 9909 39200
rect 9973 39136 9989 39200
rect 10053 39136 10069 39200
rect 10133 39136 10139 39200
rect 9823 39135 10139 39136
rect 14262 39200 14578 39201
rect 14262 39136 14268 39200
rect 14332 39136 14348 39200
rect 14412 39136 14428 39200
rect 14492 39136 14508 39200
rect 14572 39136 14578 39200
rect 14262 39135 14578 39136
rect 18701 39200 19017 39201
rect 18701 39136 18707 39200
rect 18771 39136 18787 39200
rect 18851 39136 18867 39200
rect 18931 39136 18947 39200
rect 19011 39136 19017 39200
rect 18701 39135 19017 39136
rect 3165 38656 3481 38657
rect 3165 38592 3171 38656
rect 3235 38592 3251 38656
rect 3315 38592 3331 38656
rect 3395 38592 3411 38656
rect 3475 38592 3481 38656
rect 3165 38591 3481 38592
rect 7604 38656 7920 38657
rect 7604 38592 7610 38656
rect 7674 38592 7690 38656
rect 7754 38592 7770 38656
rect 7834 38592 7850 38656
rect 7914 38592 7920 38656
rect 7604 38591 7920 38592
rect 12043 38656 12359 38657
rect 12043 38592 12049 38656
rect 12113 38592 12129 38656
rect 12193 38592 12209 38656
rect 12273 38592 12289 38656
rect 12353 38592 12359 38656
rect 12043 38591 12359 38592
rect 16482 38656 16798 38657
rect 16482 38592 16488 38656
rect 16552 38592 16568 38656
rect 16632 38592 16648 38656
rect 16712 38592 16728 38656
rect 16792 38592 16798 38656
rect 16482 38591 16798 38592
rect 5384 38112 5700 38113
rect 5384 38048 5390 38112
rect 5454 38048 5470 38112
rect 5534 38048 5550 38112
rect 5614 38048 5630 38112
rect 5694 38048 5700 38112
rect 5384 38047 5700 38048
rect 9823 38112 10139 38113
rect 9823 38048 9829 38112
rect 9893 38048 9909 38112
rect 9973 38048 9989 38112
rect 10053 38048 10069 38112
rect 10133 38048 10139 38112
rect 9823 38047 10139 38048
rect 14262 38112 14578 38113
rect 14262 38048 14268 38112
rect 14332 38048 14348 38112
rect 14412 38048 14428 38112
rect 14492 38048 14508 38112
rect 14572 38048 14578 38112
rect 14262 38047 14578 38048
rect 18701 38112 19017 38113
rect 18701 38048 18707 38112
rect 18771 38048 18787 38112
rect 18851 38048 18867 38112
rect 18931 38048 18947 38112
rect 19011 38048 19017 38112
rect 18701 38047 19017 38048
rect 3165 37568 3481 37569
rect 3165 37504 3171 37568
rect 3235 37504 3251 37568
rect 3315 37504 3331 37568
rect 3395 37504 3411 37568
rect 3475 37504 3481 37568
rect 3165 37503 3481 37504
rect 7604 37568 7920 37569
rect 7604 37504 7610 37568
rect 7674 37504 7690 37568
rect 7754 37504 7770 37568
rect 7834 37504 7850 37568
rect 7914 37504 7920 37568
rect 7604 37503 7920 37504
rect 12043 37568 12359 37569
rect 12043 37504 12049 37568
rect 12113 37504 12129 37568
rect 12193 37504 12209 37568
rect 12273 37504 12289 37568
rect 12353 37504 12359 37568
rect 12043 37503 12359 37504
rect 16482 37568 16798 37569
rect 16482 37504 16488 37568
rect 16552 37504 16568 37568
rect 16632 37504 16648 37568
rect 16712 37504 16728 37568
rect 16792 37504 16798 37568
rect 16482 37503 16798 37504
rect 5384 37024 5700 37025
rect 5384 36960 5390 37024
rect 5454 36960 5470 37024
rect 5534 36960 5550 37024
rect 5614 36960 5630 37024
rect 5694 36960 5700 37024
rect 5384 36959 5700 36960
rect 9823 37024 10139 37025
rect 9823 36960 9829 37024
rect 9893 36960 9909 37024
rect 9973 36960 9989 37024
rect 10053 36960 10069 37024
rect 10133 36960 10139 37024
rect 9823 36959 10139 36960
rect 14262 37024 14578 37025
rect 14262 36960 14268 37024
rect 14332 36960 14348 37024
rect 14412 36960 14428 37024
rect 14492 36960 14508 37024
rect 14572 36960 14578 37024
rect 14262 36959 14578 36960
rect 18701 37024 19017 37025
rect 18701 36960 18707 37024
rect 18771 36960 18787 37024
rect 18851 36960 18867 37024
rect 18931 36960 18947 37024
rect 19011 36960 19017 37024
rect 18701 36959 19017 36960
rect 3165 36480 3481 36481
rect 3165 36416 3171 36480
rect 3235 36416 3251 36480
rect 3315 36416 3331 36480
rect 3395 36416 3411 36480
rect 3475 36416 3481 36480
rect 3165 36415 3481 36416
rect 7604 36480 7920 36481
rect 7604 36416 7610 36480
rect 7674 36416 7690 36480
rect 7754 36416 7770 36480
rect 7834 36416 7850 36480
rect 7914 36416 7920 36480
rect 7604 36415 7920 36416
rect 12043 36480 12359 36481
rect 12043 36416 12049 36480
rect 12113 36416 12129 36480
rect 12193 36416 12209 36480
rect 12273 36416 12289 36480
rect 12353 36416 12359 36480
rect 12043 36415 12359 36416
rect 16482 36480 16798 36481
rect 16482 36416 16488 36480
rect 16552 36416 16568 36480
rect 16632 36416 16648 36480
rect 16712 36416 16728 36480
rect 16792 36416 16798 36480
rect 16482 36415 16798 36416
rect 5384 35936 5700 35937
rect 5384 35872 5390 35936
rect 5454 35872 5470 35936
rect 5534 35872 5550 35936
rect 5614 35872 5630 35936
rect 5694 35872 5700 35936
rect 5384 35871 5700 35872
rect 9823 35936 10139 35937
rect 9823 35872 9829 35936
rect 9893 35872 9909 35936
rect 9973 35872 9989 35936
rect 10053 35872 10069 35936
rect 10133 35872 10139 35936
rect 9823 35871 10139 35872
rect 14262 35936 14578 35937
rect 14262 35872 14268 35936
rect 14332 35872 14348 35936
rect 14412 35872 14428 35936
rect 14492 35872 14508 35936
rect 14572 35872 14578 35936
rect 14262 35871 14578 35872
rect 18701 35936 19017 35937
rect 18701 35872 18707 35936
rect 18771 35872 18787 35936
rect 18851 35872 18867 35936
rect 18931 35872 18947 35936
rect 19011 35872 19017 35936
rect 18701 35871 19017 35872
rect 3165 35392 3481 35393
rect 3165 35328 3171 35392
rect 3235 35328 3251 35392
rect 3315 35328 3331 35392
rect 3395 35328 3411 35392
rect 3475 35328 3481 35392
rect 3165 35327 3481 35328
rect 7604 35392 7920 35393
rect 7604 35328 7610 35392
rect 7674 35328 7690 35392
rect 7754 35328 7770 35392
rect 7834 35328 7850 35392
rect 7914 35328 7920 35392
rect 7604 35327 7920 35328
rect 12043 35392 12359 35393
rect 12043 35328 12049 35392
rect 12113 35328 12129 35392
rect 12193 35328 12209 35392
rect 12273 35328 12289 35392
rect 12353 35328 12359 35392
rect 12043 35327 12359 35328
rect 16482 35392 16798 35393
rect 16482 35328 16488 35392
rect 16552 35328 16568 35392
rect 16632 35328 16648 35392
rect 16712 35328 16728 35392
rect 16792 35328 16798 35392
rect 16482 35327 16798 35328
rect 5384 34848 5700 34849
rect 5384 34784 5390 34848
rect 5454 34784 5470 34848
rect 5534 34784 5550 34848
rect 5614 34784 5630 34848
rect 5694 34784 5700 34848
rect 5384 34783 5700 34784
rect 9823 34848 10139 34849
rect 9823 34784 9829 34848
rect 9893 34784 9909 34848
rect 9973 34784 9989 34848
rect 10053 34784 10069 34848
rect 10133 34784 10139 34848
rect 9823 34783 10139 34784
rect 14262 34848 14578 34849
rect 14262 34784 14268 34848
rect 14332 34784 14348 34848
rect 14412 34784 14428 34848
rect 14492 34784 14508 34848
rect 14572 34784 14578 34848
rect 14262 34783 14578 34784
rect 18701 34848 19017 34849
rect 18701 34784 18707 34848
rect 18771 34784 18787 34848
rect 18851 34784 18867 34848
rect 18931 34784 18947 34848
rect 19011 34784 19017 34848
rect 18701 34783 19017 34784
rect 18505 34370 18571 34373
rect 19200 34370 20000 34400
rect 18505 34368 20000 34370
rect 18505 34312 18510 34368
rect 18566 34312 20000 34368
rect 18505 34310 20000 34312
rect 18505 34307 18571 34310
rect 3165 34304 3481 34305
rect 3165 34240 3171 34304
rect 3235 34240 3251 34304
rect 3315 34240 3331 34304
rect 3395 34240 3411 34304
rect 3475 34240 3481 34304
rect 3165 34239 3481 34240
rect 7604 34304 7920 34305
rect 7604 34240 7610 34304
rect 7674 34240 7690 34304
rect 7754 34240 7770 34304
rect 7834 34240 7850 34304
rect 7914 34240 7920 34304
rect 7604 34239 7920 34240
rect 12043 34304 12359 34305
rect 12043 34240 12049 34304
rect 12113 34240 12129 34304
rect 12193 34240 12209 34304
rect 12273 34240 12289 34304
rect 12353 34240 12359 34304
rect 12043 34239 12359 34240
rect 16482 34304 16798 34305
rect 16482 34240 16488 34304
rect 16552 34240 16568 34304
rect 16632 34240 16648 34304
rect 16712 34240 16728 34304
rect 16792 34240 16798 34304
rect 19200 34280 20000 34310
rect 16482 34239 16798 34240
rect 5384 33760 5700 33761
rect 5384 33696 5390 33760
rect 5454 33696 5470 33760
rect 5534 33696 5550 33760
rect 5614 33696 5630 33760
rect 5694 33696 5700 33760
rect 5384 33695 5700 33696
rect 9823 33760 10139 33761
rect 9823 33696 9829 33760
rect 9893 33696 9909 33760
rect 9973 33696 9989 33760
rect 10053 33696 10069 33760
rect 10133 33696 10139 33760
rect 9823 33695 10139 33696
rect 14262 33760 14578 33761
rect 14262 33696 14268 33760
rect 14332 33696 14348 33760
rect 14412 33696 14428 33760
rect 14492 33696 14508 33760
rect 14572 33696 14578 33760
rect 14262 33695 14578 33696
rect 18701 33760 19017 33761
rect 18701 33696 18707 33760
rect 18771 33696 18787 33760
rect 18851 33696 18867 33760
rect 18931 33696 18947 33760
rect 19011 33696 19017 33760
rect 18701 33695 19017 33696
rect 3165 33216 3481 33217
rect 3165 33152 3171 33216
rect 3235 33152 3251 33216
rect 3315 33152 3331 33216
rect 3395 33152 3411 33216
rect 3475 33152 3481 33216
rect 3165 33151 3481 33152
rect 7604 33216 7920 33217
rect 7604 33152 7610 33216
rect 7674 33152 7690 33216
rect 7754 33152 7770 33216
rect 7834 33152 7850 33216
rect 7914 33152 7920 33216
rect 7604 33151 7920 33152
rect 12043 33216 12359 33217
rect 12043 33152 12049 33216
rect 12113 33152 12129 33216
rect 12193 33152 12209 33216
rect 12273 33152 12289 33216
rect 12353 33152 12359 33216
rect 12043 33151 12359 33152
rect 16482 33216 16798 33217
rect 16482 33152 16488 33216
rect 16552 33152 16568 33216
rect 16632 33152 16648 33216
rect 16712 33152 16728 33216
rect 16792 33152 16798 33216
rect 16482 33151 16798 33152
rect 5384 32672 5700 32673
rect 5384 32608 5390 32672
rect 5454 32608 5470 32672
rect 5534 32608 5550 32672
rect 5614 32608 5630 32672
rect 5694 32608 5700 32672
rect 5384 32607 5700 32608
rect 9823 32672 10139 32673
rect 9823 32608 9829 32672
rect 9893 32608 9909 32672
rect 9973 32608 9989 32672
rect 10053 32608 10069 32672
rect 10133 32608 10139 32672
rect 9823 32607 10139 32608
rect 14262 32672 14578 32673
rect 14262 32608 14268 32672
rect 14332 32608 14348 32672
rect 14412 32608 14428 32672
rect 14492 32608 14508 32672
rect 14572 32608 14578 32672
rect 14262 32607 14578 32608
rect 18701 32672 19017 32673
rect 18701 32608 18707 32672
rect 18771 32608 18787 32672
rect 18851 32608 18867 32672
rect 18931 32608 18947 32672
rect 19011 32608 19017 32672
rect 18701 32607 19017 32608
rect 3165 32128 3481 32129
rect 3165 32064 3171 32128
rect 3235 32064 3251 32128
rect 3315 32064 3331 32128
rect 3395 32064 3411 32128
rect 3475 32064 3481 32128
rect 3165 32063 3481 32064
rect 7604 32128 7920 32129
rect 7604 32064 7610 32128
rect 7674 32064 7690 32128
rect 7754 32064 7770 32128
rect 7834 32064 7850 32128
rect 7914 32064 7920 32128
rect 7604 32063 7920 32064
rect 12043 32128 12359 32129
rect 12043 32064 12049 32128
rect 12113 32064 12129 32128
rect 12193 32064 12209 32128
rect 12273 32064 12289 32128
rect 12353 32064 12359 32128
rect 12043 32063 12359 32064
rect 16482 32128 16798 32129
rect 16482 32064 16488 32128
rect 16552 32064 16568 32128
rect 16632 32064 16648 32128
rect 16712 32064 16728 32128
rect 16792 32064 16798 32128
rect 16482 32063 16798 32064
rect 5384 31584 5700 31585
rect 5384 31520 5390 31584
rect 5454 31520 5470 31584
rect 5534 31520 5550 31584
rect 5614 31520 5630 31584
rect 5694 31520 5700 31584
rect 5384 31519 5700 31520
rect 9823 31584 10139 31585
rect 9823 31520 9829 31584
rect 9893 31520 9909 31584
rect 9973 31520 9989 31584
rect 10053 31520 10069 31584
rect 10133 31520 10139 31584
rect 9823 31519 10139 31520
rect 14262 31584 14578 31585
rect 14262 31520 14268 31584
rect 14332 31520 14348 31584
rect 14412 31520 14428 31584
rect 14492 31520 14508 31584
rect 14572 31520 14578 31584
rect 14262 31519 14578 31520
rect 18701 31584 19017 31585
rect 18701 31520 18707 31584
rect 18771 31520 18787 31584
rect 18851 31520 18867 31584
rect 18931 31520 18947 31584
rect 19011 31520 19017 31584
rect 18701 31519 19017 31520
rect 3165 31040 3481 31041
rect 3165 30976 3171 31040
rect 3235 30976 3251 31040
rect 3315 30976 3331 31040
rect 3395 30976 3411 31040
rect 3475 30976 3481 31040
rect 3165 30975 3481 30976
rect 7604 31040 7920 31041
rect 7604 30976 7610 31040
rect 7674 30976 7690 31040
rect 7754 30976 7770 31040
rect 7834 30976 7850 31040
rect 7914 30976 7920 31040
rect 7604 30975 7920 30976
rect 12043 31040 12359 31041
rect 12043 30976 12049 31040
rect 12113 30976 12129 31040
rect 12193 30976 12209 31040
rect 12273 30976 12289 31040
rect 12353 30976 12359 31040
rect 12043 30975 12359 30976
rect 16482 31040 16798 31041
rect 16482 30976 16488 31040
rect 16552 30976 16568 31040
rect 16632 30976 16648 31040
rect 16712 30976 16728 31040
rect 16792 30976 16798 31040
rect 16482 30975 16798 30976
rect 5384 30496 5700 30497
rect 5384 30432 5390 30496
rect 5454 30432 5470 30496
rect 5534 30432 5550 30496
rect 5614 30432 5630 30496
rect 5694 30432 5700 30496
rect 5384 30431 5700 30432
rect 9823 30496 10139 30497
rect 9823 30432 9829 30496
rect 9893 30432 9909 30496
rect 9973 30432 9989 30496
rect 10053 30432 10069 30496
rect 10133 30432 10139 30496
rect 9823 30431 10139 30432
rect 14262 30496 14578 30497
rect 14262 30432 14268 30496
rect 14332 30432 14348 30496
rect 14412 30432 14428 30496
rect 14492 30432 14508 30496
rect 14572 30432 14578 30496
rect 14262 30431 14578 30432
rect 18701 30496 19017 30497
rect 18701 30432 18707 30496
rect 18771 30432 18787 30496
rect 18851 30432 18867 30496
rect 18931 30432 18947 30496
rect 19011 30432 19017 30496
rect 18701 30431 19017 30432
rect 3165 29952 3481 29953
rect 3165 29888 3171 29952
rect 3235 29888 3251 29952
rect 3315 29888 3331 29952
rect 3395 29888 3411 29952
rect 3475 29888 3481 29952
rect 3165 29887 3481 29888
rect 7604 29952 7920 29953
rect 7604 29888 7610 29952
rect 7674 29888 7690 29952
rect 7754 29888 7770 29952
rect 7834 29888 7850 29952
rect 7914 29888 7920 29952
rect 7604 29887 7920 29888
rect 12043 29952 12359 29953
rect 12043 29888 12049 29952
rect 12113 29888 12129 29952
rect 12193 29888 12209 29952
rect 12273 29888 12289 29952
rect 12353 29888 12359 29952
rect 12043 29887 12359 29888
rect 16482 29952 16798 29953
rect 16482 29888 16488 29952
rect 16552 29888 16568 29952
rect 16632 29888 16648 29952
rect 16712 29888 16728 29952
rect 16792 29888 16798 29952
rect 16482 29887 16798 29888
rect 5384 29408 5700 29409
rect 5384 29344 5390 29408
rect 5454 29344 5470 29408
rect 5534 29344 5550 29408
rect 5614 29344 5630 29408
rect 5694 29344 5700 29408
rect 5384 29343 5700 29344
rect 9823 29408 10139 29409
rect 9823 29344 9829 29408
rect 9893 29344 9909 29408
rect 9973 29344 9989 29408
rect 10053 29344 10069 29408
rect 10133 29344 10139 29408
rect 9823 29343 10139 29344
rect 14262 29408 14578 29409
rect 14262 29344 14268 29408
rect 14332 29344 14348 29408
rect 14412 29344 14428 29408
rect 14492 29344 14508 29408
rect 14572 29344 14578 29408
rect 14262 29343 14578 29344
rect 18701 29408 19017 29409
rect 18701 29344 18707 29408
rect 18771 29344 18787 29408
rect 18851 29344 18867 29408
rect 18931 29344 18947 29408
rect 19011 29344 19017 29408
rect 18701 29343 19017 29344
rect 3165 28864 3481 28865
rect 3165 28800 3171 28864
rect 3235 28800 3251 28864
rect 3315 28800 3331 28864
rect 3395 28800 3411 28864
rect 3475 28800 3481 28864
rect 3165 28799 3481 28800
rect 7604 28864 7920 28865
rect 7604 28800 7610 28864
rect 7674 28800 7690 28864
rect 7754 28800 7770 28864
rect 7834 28800 7850 28864
rect 7914 28800 7920 28864
rect 7604 28799 7920 28800
rect 12043 28864 12359 28865
rect 12043 28800 12049 28864
rect 12113 28800 12129 28864
rect 12193 28800 12209 28864
rect 12273 28800 12289 28864
rect 12353 28800 12359 28864
rect 12043 28799 12359 28800
rect 16482 28864 16798 28865
rect 16482 28800 16488 28864
rect 16552 28800 16568 28864
rect 16632 28800 16648 28864
rect 16712 28800 16728 28864
rect 16792 28800 16798 28864
rect 16482 28799 16798 28800
rect 5384 28320 5700 28321
rect 5384 28256 5390 28320
rect 5454 28256 5470 28320
rect 5534 28256 5550 28320
rect 5614 28256 5630 28320
rect 5694 28256 5700 28320
rect 5384 28255 5700 28256
rect 9823 28320 10139 28321
rect 9823 28256 9829 28320
rect 9893 28256 9909 28320
rect 9973 28256 9989 28320
rect 10053 28256 10069 28320
rect 10133 28256 10139 28320
rect 9823 28255 10139 28256
rect 14262 28320 14578 28321
rect 14262 28256 14268 28320
rect 14332 28256 14348 28320
rect 14412 28256 14428 28320
rect 14492 28256 14508 28320
rect 14572 28256 14578 28320
rect 14262 28255 14578 28256
rect 18701 28320 19017 28321
rect 18701 28256 18707 28320
rect 18771 28256 18787 28320
rect 18851 28256 18867 28320
rect 18931 28256 18947 28320
rect 19011 28256 19017 28320
rect 18701 28255 19017 28256
rect 18597 28114 18663 28117
rect 19200 28114 20000 28144
rect 18597 28112 20000 28114
rect 18597 28056 18602 28112
rect 18658 28056 20000 28112
rect 18597 28054 20000 28056
rect 18597 28051 18663 28054
rect 19200 28024 20000 28054
rect 3165 27776 3481 27777
rect 3165 27712 3171 27776
rect 3235 27712 3251 27776
rect 3315 27712 3331 27776
rect 3395 27712 3411 27776
rect 3475 27712 3481 27776
rect 3165 27711 3481 27712
rect 7604 27776 7920 27777
rect 7604 27712 7610 27776
rect 7674 27712 7690 27776
rect 7754 27712 7770 27776
rect 7834 27712 7850 27776
rect 7914 27712 7920 27776
rect 7604 27711 7920 27712
rect 12043 27776 12359 27777
rect 12043 27712 12049 27776
rect 12113 27712 12129 27776
rect 12193 27712 12209 27776
rect 12273 27712 12289 27776
rect 12353 27712 12359 27776
rect 12043 27711 12359 27712
rect 16482 27776 16798 27777
rect 16482 27712 16488 27776
rect 16552 27712 16568 27776
rect 16632 27712 16648 27776
rect 16712 27712 16728 27776
rect 16792 27712 16798 27776
rect 16482 27711 16798 27712
rect 5384 27232 5700 27233
rect 5384 27168 5390 27232
rect 5454 27168 5470 27232
rect 5534 27168 5550 27232
rect 5614 27168 5630 27232
rect 5694 27168 5700 27232
rect 5384 27167 5700 27168
rect 9823 27232 10139 27233
rect 9823 27168 9829 27232
rect 9893 27168 9909 27232
rect 9973 27168 9989 27232
rect 10053 27168 10069 27232
rect 10133 27168 10139 27232
rect 9823 27167 10139 27168
rect 14262 27232 14578 27233
rect 14262 27168 14268 27232
rect 14332 27168 14348 27232
rect 14412 27168 14428 27232
rect 14492 27168 14508 27232
rect 14572 27168 14578 27232
rect 14262 27167 14578 27168
rect 18701 27232 19017 27233
rect 18701 27168 18707 27232
rect 18771 27168 18787 27232
rect 18851 27168 18867 27232
rect 18931 27168 18947 27232
rect 19011 27168 19017 27232
rect 18701 27167 19017 27168
rect 3165 26688 3481 26689
rect 3165 26624 3171 26688
rect 3235 26624 3251 26688
rect 3315 26624 3331 26688
rect 3395 26624 3411 26688
rect 3475 26624 3481 26688
rect 3165 26623 3481 26624
rect 7604 26688 7920 26689
rect 7604 26624 7610 26688
rect 7674 26624 7690 26688
rect 7754 26624 7770 26688
rect 7834 26624 7850 26688
rect 7914 26624 7920 26688
rect 7604 26623 7920 26624
rect 12043 26688 12359 26689
rect 12043 26624 12049 26688
rect 12113 26624 12129 26688
rect 12193 26624 12209 26688
rect 12273 26624 12289 26688
rect 12353 26624 12359 26688
rect 12043 26623 12359 26624
rect 16482 26688 16798 26689
rect 16482 26624 16488 26688
rect 16552 26624 16568 26688
rect 16632 26624 16648 26688
rect 16712 26624 16728 26688
rect 16792 26624 16798 26688
rect 16482 26623 16798 26624
rect 5384 26144 5700 26145
rect 5384 26080 5390 26144
rect 5454 26080 5470 26144
rect 5534 26080 5550 26144
rect 5614 26080 5630 26144
rect 5694 26080 5700 26144
rect 5384 26079 5700 26080
rect 9823 26144 10139 26145
rect 9823 26080 9829 26144
rect 9893 26080 9909 26144
rect 9973 26080 9989 26144
rect 10053 26080 10069 26144
rect 10133 26080 10139 26144
rect 9823 26079 10139 26080
rect 14262 26144 14578 26145
rect 14262 26080 14268 26144
rect 14332 26080 14348 26144
rect 14412 26080 14428 26144
rect 14492 26080 14508 26144
rect 14572 26080 14578 26144
rect 14262 26079 14578 26080
rect 18701 26144 19017 26145
rect 18701 26080 18707 26144
rect 18771 26080 18787 26144
rect 18851 26080 18867 26144
rect 18931 26080 18947 26144
rect 19011 26080 19017 26144
rect 18701 26079 19017 26080
rect 3165 25600 3481 25601
rect 3165 25536 3171 25600
rect 3235 25536 3251 25600
rect 3315 25536 3331 25600
rect 3395 25536 3411 25600
rect 3475 25536 3481 25600
rect 3165 25535 3481 25536
rect 7604 25600 7920 25601
rect 7604 25536 7610 25600
rect 7674 25536 7690 25600
rect 7754 25536 7770 25600
rect 7834 25536 7850 25600
rect 7914 25536 7920 25600
rect 7604 25535 7920 25536
rect 12043 25600 12359 25601
rect 12043 25536 12049 25600
rect 12113 25536 12129 25600
rect 12193 25536 12209 25600
rect 12273 25536 12289 25600
rect 12353 25536 12359 25600
rect 12043 25535 12359 25536
rect 16482 25600 16798 25601
rect 16482 25536 16488 25600
rect 16552 25536 16568 25600
rect 16632 25536 16648 25600
rect 16712 25536 16728 25600
rect 16792 25536 16798 25600
rect 16482 25535 16798 25536
rect 5384 25056 5700 25057
rect 5384 24992 5390 25056
rect 5454 24992 5470 25056
rect 5534 24992 5550 25056
rect 5614 24992 5630 25056
rect 5694 24992 5700 25056
rect 5384 24991 5700 24992
rect 9823 25056 10139 25057
rect 9823 24992 9829 25056
rect 9893 24992 9909 25056
rect 9973 24992 9989 25056
rect 10053 24992 10069 25056
rect 10133 24992 10139 25056
rect 9823 24991 10139 24992
rect 14262 25056 14578 25057
rect 14262 24992 14268 25056
rect 14332 24992 14348 25056
rect 14412 24992 14428 25056
rect 14492 24992 14508 25056
rect 14572 24992 14578 25056
rect 14262 24991 14578 24992
rect 18701 25056 19017 25057
rect 18701 24992 18707 25056
rect 18771 24992 18787 25056
rect 18851 24992 18867 25056
rect 18931 24992 18947 25056
rect 19011 24992 19017 25056
rect 18701 24991 19017 24992
rect 3165 24512 3481 24513
rect 3165 24448 3171 24512
rect 3235 24448 3251 24512
rect 3315 24448 3331 24512
rect 3395 24448 3411 24512
rect 3475 24448 3481 24512
rect 3165 24447 3481 24448
rect 7604 24512 7920 24513
rect 7604 24448 7610 24512
rect 7674 24448 7690 24512
rect 7754 24448 7770 24512
rect 7834 24448 7850 24512
rect 7914 24448 7920 24512
rect 7604 24447 7920 24448
rect 12043 24512 12359 24513
rect 12043 24448 12049 24512
rect 12113 24448 12129 24512
rect 12193 24448 12209 24512
rect 12273 24448 12289 24512
rect 12353 24448 12359 24512
rect 12043 24447 12359 24448
rect 16482 24512 16798 24513
rect 16482 24448 16488 24512
rect 16552 24448 16568 24512
rect 16632 24448 16648 24512
rect 16712 24448 16728 24512
rect 16792 24448 16798 24512
rect 16482 24447 16798 24448
rect 5384 23968 5700 23969
rect 5384 23904 5390 23968
rect 5454 23904 5470 23968
rect 5534 23904 5550 23968
rect 5614 23904 5630 23968
rect 5694 23904 5700 23968
rect 5384 23903 5700 23904
rect 9823 23968 10139 23969
rect 9823 23904 9829 23968
rect 9893 23904 9909 23968
rect 9973 23904 9989 23968
rect 10053 23904 10069 23968
rect 10133 23904 10139 23968
rect 9823 23903 10139 23904
rect 14262 23968 14578 23969
rect 14262 23904 14268 23968
rect 14332 23904 14348 23968
rect 14412 23904 14428 23968
rect 14492 23904 14508 23968
rect 14572 23904 14578 23968
rect 14262 23903 14578 23904
rect 18701 23968 19017 23969
rect 18701 23904 18707 23968
rect 18771 23904 18787 23968
rect 18851 23904 18867 23968
rect 18931 23904 18947 23968
rect 19011 23904 19017 23968
rect 18701 23903 19017 23904
rect 3165 23424 3481 23425
rect 3165 23360 3171 23424
rect 3235 23360 3251 23424
rect 3315 23360 3331 23424
rect 3395 23360 3411 23424
rect 3475 23360 3481 23424
rect 3165 23359 3481 23360
rect 7604 23424 7920 23425
rect 7604 23360 7610 23424
rect 7674 23360 7690 23424
rect 7754 23360 7770 23424
rect 7834 23360 7850 23424
rect 7914 23360 7920 23424
rect 7604 23359 7920 23360
rect 12043 23424 12359 23425
rect 12043 23360 12049 23424
rect 12113 23360 12129 23424
rect 12193 23360 12209 23424
rect 12273 23360 12289 23424
rect 12353 23360 12359 23424
rect 12043 23359 12359 23360
rect 16482 23424 16798 23425
rect 16482 23360 16488 23424
rect 16552 23360 16568 23424
rect 16632 23360 16648 23424
rect 16712 23360 16728 23424
rect 16792 23360 16798 23424
rect 16482 23359 16798 23360
rect 5384 22880 5700 22881
rect 5384 22816 5390 22880
rect 5454 22816 5470 22880
rect 5534 22816 5550 22880
rect 5614 22816 5630 22880
rect 5694 22816 5700 22880
rect 5384 22815 5700 22816
rect 9823 22880 10139 22881
rect 9823 22816 9829 22880
rect 9893 22816 9909 22880
rect 9973 22816 9989 22880
rect 10053 22816 10069 22880
rect 10133 22816 10139 22880
rect 9823 22815 10139 22816
rect 14262 22880 14578 22881
rect 14262 22816 14268 22880
rect 14332 22816 14348 22880
rect 14412 22816 14428 22880
rect 14492 22816 14508 22880
rect 14572 22816 14578 22880
rect 14262 22815 14578 22816
rect 18701 22880 19017 22881
rect 18701 22816 18707 22880
rect 18771 22816 18787 22880
rect 18851 22816 18867 22880
rect 18931 22816 18947 22880
rect 19011 22816 19017 22880
rect 18701 22815 19017 22816
rect 3165 22336 3481 22337
rect 3165 22272 3171 22336
rect 3235 22272 3251 22336
rect 3315 22272 3331 22336
rect 3395 22272 3411 22336
rect 3475 22272 3481 22336
rect 3165 22271 3481 22272
rect 7604 22336 7920 22337
rect 7604 22272 7610 22336
rect 7674 22272 7690 22336
rect 7754 22272 7770 22336
rect 7834 22272 7850 22336
rect 7914 22272 7920 22336
rect 7604 22271 7920 22272
rect 12043 22336 12359 22337
rect 12043 22272 12049 22336
rect 12113 22272 12129 22336
rect 12193 22272 12209 22336
rect 12273 22272 12289 22336
rect 12353 22272 12359 22336
rect 12043 22271 12359 22272
rect 16482 22336 16798 22337
rect 16482 22272 16488 22336
rect 16552 22272 16568 22336
rect 16632 22272 16648 22336
rect 16712 22272 16728 22336
rect 16792 22272 16798 22336
rect 16482 22271 16798 22272
rect 18505 22130 18571 22133
rect 18505 22128 19626 22130
rect 18505 22072 18510 22128
rect 18566 22072 19626 22128
rect 18505 22070 19626 22072
rect 18505 22067 18571 22070
rect 19566 21888 19626 22070
rect 5384 21792 5700 21793
rect 5384 21728 5390 21792
rect 5454 21728 5470 21792
rect 5534 21728 5550 21792
rect 5614 21728 5630 21792
rect 5694 21728 5700 21792
rect 5384 21727 5700 21728
rect 9823 21792 10139 21793
rect 9823 21728 9829 21792
rect 9893 21728 9909 21792
rect 9973 21728 9989 21792
rect 10053 21728 10069 21792
rect 10133 21728 10139 21792
rect 9823 21727 10139 21728
rect 14262 21792 14578 21793
rect 14262 21728 14268 21792
rect 14332 21728 14348 21792
rect 14412 21728 14428 21792
rect 14492 21728 14508 21792
rect 14572 21728 14578 21792
rect 14262 21727 14578 21728
rect 18701 21792 19017 21793
rect 18701 21728 18707 21792
rect 18771 21728 18787 21792
rect 18851 21728 18867 21792
rect 18931 21728 18947 21792
rect 19011 21728 19017 21792
rect 19200 21768 20000 21888
rect 18701 21727 19017 21728
rect 3165 21248 3481 21249
rect 3165 21184 3171 21248
rect 3235 21184 3251 21248
rect 3315 21184 3331 21248
rect 3395 21184 3411 21248
rect 3475 21184 3481 21248
rect 3165 21183 3481 21184
rect 7604 21248 7920 21249
rect 7604 21184 7610 21248
rect 7674 21184 7690 21248
rect 7754 21184 7770 21248
rect 7834 21184 7850 21248
rect 7914 21184 7920 21248
rect 7604 21183 7920 21184
rect 12043 21248 12359 21249
rect 12043 21184 12049 21248
rect 12113 21184 12129 21248
rect 12193 21184 12209 21248
rect 12273 21184 12289 21248
rect 12353 21184 12359 21248
rect 12043 21183 12359 21184
rect 16482 21248 16798 21249
rect 16482 21184 16488 21248
rect 16552 21184 16568 21248
rect 16632 21184 16648 21248
rect 16712 21184 16728 21248
rect 16792 21184 16798 21248
rect 16482 21183 16798 21184
rect 5384 20704 5700 20705
rect 5384 20640 5390 20704
rect 5454 20640 5470 20704
rect 5534 20640 5550 20704
rect 5614 20640 5630 20704
rect 5694 20640 5700 20704
rect 5384 20639 5700 20640
rect 9823 20704 10139 20705
rect 9823 20640 9829 20704
rect 9893 20640 9909 20704
rect 9973 20640 9989 20704
rect 10053 20640 10069 20704
rect 10133 20640 10139 20704
rect 9823 20639 10139 20640
rect 14262 20704 14578 20705
rect 14262 20640 14268 20704
rect 14332 20640 14348 20704
rect 14412 20640 14428 20704
rect 14492 20640 14508 20704
rect 14572 20640 14578 20704
rect 14262 20639 14578 20640
rect 18701 20704 19017 20705
rect 18701 20640 18707 20704
rect 18771 20640 18787 20704
rect 18851 20640 18867 20704
rect 18931 20640 18947 20704
rect 19011 20640 19017 20704
rect 18701 20639 19017 20640
rect 3165 20160 3481 20161
rect 3165 20096 3171 20160
rect 3235 20096 3251 20160
rect 3315 20096 3331 20160
rect 3395 20096 3411 20160
rect 3475 20096 3481 20160
rect 3165 20095 3481 20096
rect 7604 20160 7920 20161
rect 7604 20096 7610 20160
rect 7674 20096 7690 20160
rect 7754 20096 7770 20160
rect 7834 20096 7850 20160
rect 7914 20096 7920 20160
rect 7604 20095 7920 20096
rect 12043 20160 12359 20161
rect 12043 20096 12049 20160
rect 12113 20096 12129 20160
rect 12193 20096 12209 20160
rect 12273 20096 12289 20160
rect 12353 20096 12359 20160
rect 12043 20095 12359 20096
rect 16482 20160 16798 20161
rect 16482 20096 16488 20160
rect 16552 20096 16568 20160
rect 16632 20096 16648 20160
rect 16712 20096 16728 20160
rect 16792 20096 16798 20160
rect 16482 20095 16798 20096
rect 5384 19616 5700 19617
rect 5384 19552 5390 19616
rect 5454 19552 5470 19616
rect 5534 19552 5550 19616
rect 5614 19552 5630 19616
rect 5694 19552 5700 19616
rect 5384 19551 5700 19552
rect 9823 19616 10139 19617
rect 9823 19552 9829 19616
rect 9893 19552 9909 19616
rect 9973 19552 9989 19616
rect 10053 19552 10069 19616
rect 10133 19552 10139 19616
rect 9823 19551 10139 19552
rect 14262 19616 14578 19617
rect 14262 19552 14268 19616
rect 14332 19552 14348 19616
rect 14412 19552 14428 19616
rect 14492 19552 14508 19616
rect 14572 19552 14578 19616
rect 14262 19551 14578 19552
rect 18701 19616 19017 19617
rect 18701 19552 18707 19616
rect 18771 19552 18787 19616
rect 18851 19552 18867 19616
rect 18931 19552 18947 19616
rect 19011 19552 19017 19616
rect 18701 19551 19017 19552
rect 3165 19072 3481 19073
rect 3165 19008 3171 19072
rect 3235 19008 3251 19072
rect 3315 19008 3331 19072
rect 3395 19008 3411 19072
rect 3475 19008 3481 19072
rect 3165 19007 3481 19008
rect 7604 19072 7920 19073
rect 7604 19008 7610 19072
rect 7674 19008 7690 19072
rect 7754 19008 7770 19072
rect 7834 19008 7850 19072
rect 7914 19008 7920 19072
rect 7604 19007 7920 19008
rect 12043 19072 12359 19073
rect 12043 19008 12049 19072
rect 12113 19008 12129 19072
rect 12193 19008 12209 19072
rect 12273 19008 12289 19072
rect 12353 19008 12359 19072
rect 12043 19007 12359 19008
rect 16482 19072 16798 19073
rect 16482 19008 16488 19072
rect 16552 19008 16568 19072
rect 16632 19008 16648 19072
rect 16712 19008 16728 19072
rect 16792 19008 16798 19072
rect 16482 19007 16798 19008
rect 5384 18528 5700 18529
rect 5384 18464 5390 18528
rect 5454 18464 5470 18528
rect 5534 18464 5550 18528
rect 5614 18464 5630 18528
rect 5694 18464 5700 18528
rect 5384 18463 5700 18464
rect 9823 18528 10139 18529
rect 9823 18464 9829 18528
rect 9893 18464 9909 18528
rect 9973 18464 9989 18528
rect 10053 18464 10069 18528
rect 10133 18464 10139 18528
rect 9823 18463 10139 18464
rect 14262 18528 14578 18529
rect 14262 18464 14268 18528
rect 14332 18464 14348 18528
rect 14412 18464 14428 18528
rect 14492 18464 14508 18528
rect 14572 18464 14578 18528
rect 14262 18463 14578 18464
rect 18701 18528 19017 18529
rect 18701 18464 18707 18528
rect 18771 18464 18787 18528
rect 18851 18464 18867 18528
rect 18931 18464 18947 18528
rect 19011 18464 19017 18528
rect 18701 18463 19017 18464
rect 3165 17984 3481 17985
rect 3165 17920 3171 17984
rect 3235 17920 3251 17984
rect 3315 17920 3331 17984
rect 3395 17920 3411 17984
rect 3475 17920 3481 17984
rect 3165 17919 3481 17920
rect 7604 17984 7920 17985
rect 7604 17920 7610 17984
rect 7674 17920 7690 17984
rect 7754 17920 7770 17984
rect 7834 17920 7850 17984
rect 7914 17920 7920 17984
rect 7604 17919 7920 17920
rect 12043 17984 12359 17985
rect 12043 17920 12049 17984
rect 12113 17920 12129 17984
rect 12193 17920 12209 17984
rect 12273 17920 12289 17984
rect 12353 17920 12359 17984
rect 12043 17919 12359 17920
rect 16482 17984 16798 17985
rect 16482 17920 16488 17984
rect 16552 17920 16568 17984
rect 16632 17920 16648 17984
rect 16712 17920 16728 17984
rect 16792 17920 16798 17984
rect 16482 17919 16798 17920
rect 5384 17440 5700 17441
rect 5384 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5700 17440
rect 5384 17375 5700 17376
rect 9823 17440 10139 17441
rect 9823 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10139 17440
rect 9823 17375 10139 17376
rect 14262 17440 14578 17441
rect 14262 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14578 17440
rect 14262 17375 14578 17376
rect 18701 17440 19017 17441
rect 18701 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19017 17440
rect 18701 17375 19017 17376
rect 3165 16896 3481 16897
rect 3165 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3481 16896
rect 3165 16831 3481 16832
rect 7604 16896 7920 16897
rect 7604 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7920 16896
rect 7604 16831 7920 16832
rect 12043 16896 12359 16897
rect 12043 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12359 16896
rect 12043 16831 12359 16832
rect 16482 16896 16798 16897
rect 16482 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16798 16896
rect 16482 16831 16798 16832
rect 5384 16352 5700 16353
rect 5384 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5700 16352
rect 5384 16287 5700 16288
rect 9823 16352 10139 16353
rect 9823 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10139 16352
rect 9823 16287 10139 16288
rect 14262 16352 14578 16353
rect 14262 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14578 16352
rect 14262 16287 14578 16288
rect 18701 16352 19017 16353
rect 18701 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19017 16352
rect 18701 16287 19017 16288
rect 3165 15808 3481 15809
rect 3165 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3481 15808
rect 3165 15743 3481 15744
rect 7604 15808 7920 15809
rect 7604 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7920 15808
rect 7604 15743 7920 15744
rect 12043 15808 12359 15809
rect 12043 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12359 15808
rect 12043 15743 12359 15744
rect 16482 15808 16798 15809
rect 16482 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16798 15808
rect 16482 15743 16798 15744
rect 18321 15602 18387 15605
rect 19200 15602 20000 15632
rect 18321 15600 20000 15602
rect 18321 15544 18326 15600
rect 18382 15544 20000 15600
rect 18321 15542 20000 15544
rect 18321 15539 18387 15542
rect 19200 15512 20000 15542
rect 5384 15264 5700 15265
rect 5384 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5700 15264
rect 5384 15199 5700 15200
rect 9823 15264 10139 15265
rect 9823 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10139 15264
rect 9823 15199 10139 15200
rect 14262 15264 14578 15265
rect 14262 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14578 15264
rect 14262 15199 14578 15200
rect 18701 15264 19017 15265
rect 18701 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19017 15264
rect 18701 15199 19017 15200
rect 3165 14720 3481 14721
rect 3165 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3481 14720
rect 3165 14655 3481 14656
rect 7604 14720 7920 14721
rect 7604 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7920 14720
rect 7604 14655 7920 14656
rect 12043 14720 12359 14721
rect 12043 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12359 14720
rect 12043 14655 12359 14656
rect 16482 14720 16798 14721
rect 16482 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16798 14720
rect 16482 14655 16798 14656
rect 5384 14176 5700 14177
rect 5384 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5700 14176
rect 5384 14111 5700 14112
rect 9823 14176 10139 14177
rect 9823 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10139 14176
rect 9823 14111 10139 14112
rect 14262 14176 14578 14177
rect 14262 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14578 14176
rect 14262 14111 14578 14112
rect 18701 14176 19017 14177
rect 18701 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19017 14176
rect 18701 14111 19017 14112
rect 3165 13632 3481 13633
rect 3165 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3481 13632
rect 3165 13567 3481 13568
rect 7604 13632 7920 13633
rect 7604 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7920 13632
rect 7604 13567 7920 13568
rect 12043 13632 12359 13633
rect 12043 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12359 13632
rect 12043 13567 12359 13568
rect 16482 13632 16798 13633
rect 16482 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16798 13632
rect 16482 13567 16798 13568
rect 5384 13088 5700 13089
rect 5384 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5700 13088
rect 5384 13023 5700 13024
rect 9823 13088 10139 13089
rect 9823 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10139 13088
rect 9823 13023 10139 13024
rect 14262 13088 14578 13089
rect 14262 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14578 13088
rect 14262 13023 14578 13024
rect 18701 13088 19017 13089
rect 18701 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19017 13088
rect 18701 13023 19017 13024
rect 3165 12544 3481 12545
rect 3165 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3481 12544
rect 3165 12479 3481 12480
rect 7604 12544 7920 12545
rect 7604 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7920 12544
rect 7604 12479 7920 12480
rect 12043 12544 12359 12545
rect 12043 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12359 12544
rect 12043 12479 12359 12480
rect 16482 12544 16798 12545
rect 16482 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16798 12544
rect 16482 12479 16798 12480
rect 5384 12000 5700 12001
rect 5384 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5700 12000
rect 5384 11935 5700 11936
rect 9823 12000 10139 12001
rect 9823 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10139 12000
rect 9823 11935 10139 11936
rect 14262 12000 14578 12001
rect 14262 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14578 12000
rect 14262 11935 14578 11936
rect 18701 12000 19017 12001
rect 18701 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19017 12000
rect 18701 11935 19017 11936
rect 3165 11456 3481 11457
rect 3165 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3481 11456
rect 3165 11391 3481 11392
rect 7604 11456 7920 11457
rect 7604 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7920 11456
rect 7604 11391 7920 11392
rect 12043 11456 12359 11457
rect 12043 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12359 11456
rect 12043 11391 12359 11392
rect 16482 11456 16798 11457
rect 16482 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16798 11456
rect 16482 11391 16798 11392
rect 5384 10912 5700 10913
rect 5384 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5700 10912
rect 5384 10847 5700 10848
rect 9823 10912 10139 10913
rect 9823 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10139 10912
rect 9823 10847 10139 10848
rect 14262 10912 14578 10913
rect 14262 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14578 10912
rect 14262 10847 14578 10848
rect 18701 10912 19017 10913
rect 18701 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19017 10912
rect 18701 10847 19017 10848
rect 3165 10368 3481 10369
rect 3165 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3481 10368
rect 3165 10303 3481 10304
rect 7604 10368 7920 10369
rect 7604 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7920 10368
rect 7604 10303 7920 10304
rect 12043 10368 12359 10369
rect 12043 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12359 10368
rect 12043 10303 12359 10304
rect 16482 10368 16798 10369
rect 16482 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16798 10368
rect 16482 10303 16798 10304
rect 5384 9824 5700 9825
rect 5384 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5700 9824
rect 5384 9759 5700 9760
rect 9823 9824 10139 9825
rect 9823 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10139 9824
rect 9823 9759 10139 9760
rect 14262 9824 14578 9825
rect 14262 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14578 9824
rect 14262 9759 14578 9760
rect 18701 9824 19017 9825
rect 18701 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19017 9824
rect 18701 9759 19017 9760
rect 18505 9346 18571 9349
rect 19200 9346 20000 9376
rect 18505 9344 20000 9346
rect 18505 9288 18510 9344
rect 18566 9288 20000 9344
rect 18505 9286 20000 9288
rect 18505 9283 18571 9286
rect 3165 9280 3481 9281
rect 3165 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3481 9280
rect 3165 9215 3481 9216
rect 7604 9280 7920 9281
rect 7604 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7920 9280
rect 7604 9215 7920 9216
rect 12043 9280 12359 9281
rect 12043 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12359 9280
rect 12043 9215 12359 9216
rect 16482 9280 16798 9281
rect 16482 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16798 9280
rect 19200 9256 20000 9286
rect 16482 9215 16798 9216
rect 5384 8736 5700 8737
rect 5384 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5700 8736
rect 5384 8671 5700 8672
rect 9823 8736 10139 8737
rect 9823 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10139 8736
rect 9823 8671 10139 8672
rect 14262 8736 14578 8737
rect 14262 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14578 8736
rect 14262 8671 14578 8672
rect 18701 8736 19017 8737
rect 18701 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19017 8736
rect 18701 8671 19017 8672
rect 3165 8192 3481 8193
rect 3165 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3481 8192
rect 3165 8127 3481 8128
rect 7604 8192 7920 8193
rect 7604 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7920 8192
rect 7604 8127 7920 8128
rect 12043 8192 12359 8193
rect 12043 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12359 8192
rect 12043 8127 12359 8128
rect 16482 8192 16798 8193
rect 16482 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16798 8192
rect 16482 8127 16798 8128
rect 5384 7648 5700 7649
rect 5384 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5700 7648
rect 5384 7583 5700 7584
rect 9823 7648 10139 7649
rect 9823 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10139 7648
rect 9823 7583 10139 7584
rect 14262 7648 14578 7649
rect 14262 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14578 7648
rect 14262 7583 14578 7584
rect 18701 7648 19017 7649
rect 18701 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19017 7648
rect 18701 7583 19017 7584
rect 3165 7104 3481 7105
rect 3165 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3481 7104
rect 3165 7039 3481 7040
rect 7604 7104 7920 7105
rect 7604 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7920 7104
rect 7604 7039 7920 7040
rect 12043 7104 12359 7105
rect 12043 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12359 7104
rect 12043 7039 12359 7040
rect 16482 7104 16798 7105
rect 16482 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16798 7104
rect 16482 7039 16798 7040
rect 5384 6560 5700 6561
rect 5384 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5700 6560
rect 5384 6495 5700 6496
rect 9823 6560 10139 6561
rect 9823 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10139 6560
rect 9823 6495 10139 6496
rect 14262 6560 14578 6561
rect 14262 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14578 6560
rect 14262 6495 14578 6496
rect 18701 6560 19017 6561
rect 18701 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19017 6560
rect 18701 6495 19017 6496
rect 3165 6016 3481 6017
rect 3165 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3481 6016
rect 3165 5951 3481 5952
rect 7604 6016 7920 6017
rect 7604 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7920 6016
rect 7604 5951 7920 5952
rect 12043 6016 12359 6017
rect 12043 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12359 6016
rect 12043 5951 12359 5952
rect 16482 6016 16798 6017
rect 16482 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16798 6016
rect 16482 5951 16798 5952
rect 5384 5472 5700 5473
rect 5384 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5700 5472
rect 5384 5407 5700 5408
rect 9823 5472 10139 5473
rect 9823 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10139 5472
rect 9823 5407 10139 5408
rect 14262 5472 14578 5473
rect 14262 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14578 5472
rect 14262 5407 14578 5408
rect 18701 5472 19017 5473
rect 18701 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19017 5472
rect 18701 5407 19017 5408
rect 3165 4928 3481 4929
rect 3165 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3481 4928
rect 3165 4863 3481 4864
rect 7604 4928 7920 4929
rect 7604 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7920 4928
rect 7604 4863 7920 4864
rect 12043 4928 12359 4929
rect 12043 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12359 4928
rect 12043 4863 12359 4864
rect 16482 4928 16798 4929
rect 16482 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16798 4928
rect 16482 4863 16798 4864
rect 5384 4384 5700 4385
rect 5384 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5700 4384
rect 5384 4319 5700 4320
rect 9823 4384 10139 4385
rect 9823 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10139 4384
rect 9823 4319 10139 4320
rect 14262 4384 14578 4385
rect 14262 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14578 4384
rect 14262 4319 14578 4320
rect 18701 4384 19017 4385
rect 18701 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19017 4384
rect 18701 4319 19017 4320
rect 3165 3840 3481 3841
rect 3165 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3481 3840
rect 3165 3775 3481 3776
rect 7604 3840 7920 3841
rect 7604 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7920 3840
rect 7604 3775 7920 3776
rect 12043 3840 12359 3841
rect 12043 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12359 3840
rect 12043 3775 12359 3776
rect 16482 3840 16798 3841
rect 16482 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16798 3840
rect 16482 3775 16798 3776
rect 5384 3296 5700 3297
rect 5384 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5700 3296
rect 5384 3231 5700 3232
rect 9823 3296 10139 3297
rect 9823 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10139 3296
rect 9823 3231 10139 3232
rect 14262 3296 14578 3297
rect 14262 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14578 3296
rect 14262 3231 14578 3232
rect 18701 3296 19017 3297
rect 18701 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19017 3296
rect 18701 3231 19017 3232
rect 18321 3090 18387 3093
rect 19200 3090 20000 3120
rect 18321 3088 20000 3090
rect 18321 3032 18326 3088
rect 18382 3032 20000 3088
rect 18321 3030 20000 3032
rect 18321 3027 18387 3030
rect 19200 3000 20000 3030
rect 3165 2752 3481 2753
rect 3165 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3481 2752
rect 3165 2687 3481 2688
rect 7604 2752 7920 2753
rect 7604 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7920 2752
rect 7604 2687 7920 2688
rect 12043 2752 12359 2753
rect 12043 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12359 2752
rect 12043 2687 12359 2688
rect 16482 2752 16798 2753
rect 16482 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16798 2752
rect 16482 2687 16798 2688
rect 5384 2208 5700 2209
rect 5384 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5700 2208
rect 5384 2143 5700 2144
rect 9823 2208 10139 2209
rect 9823 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10139 2208
rect 9823 2143 10139 2144
rect 14262 2208 14578 2209
rect 14262 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14578 2208
rect 14262 2143 14578 2144
rect 18701 2208 19017 2209
rect 18701 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19017 2208
rect 18701 2143 19017 2144
<< via3 >>
rect 3171 47356 3235 47360
rect 3171 47300 3175 47356
rect 3175 47300 3231 47356
rect 3231 47300 3235 47356
rect 3171 47296 3235 47300
rect 3251 47356 3315 47360
rect 3251 47300 3255 47356
rect 3255 47300 3311 47356
rect 3311 47300 3315 47356
rect 3251 47296 3315 47300
rect 3331 47356 3395 47360
rect 3331 47300 3335 47356
rect 3335 47300 3391 47356
rect 3391 47300 3395 47356
rect 3331 47296 3395 47300
rect 3411 47356 3475 47360
rect 3411 47300 3415 47356
rect 3415 47300 3471 47356
rect 3471 47300 3475 47356
rect 3411 47296 3475 47300
rect 7610 47356 7674 47360
rect 7610 47300 7614 47356
rect 7614 47300 7670 47356
rect 7670 47300 7674 47356
rect 7610 47296 7674 47300
rect 7690 47356 7754 47360
rect 7690 47300 7694 47356
rect 7694 47300 7750 47356
rect 7750 47300 7754 47356
rect 7690 47296 7754 47300
rect 7770 47356 7834 47360
rect 7770 47300 7774 47356
rect 7774 47300 7830 47356
rect 7830 47300 7834 47356
rect 7770 47296 7834 47300
rect 7850 47356 7914 47360
rect 7850 47300 7854 47356
rect 7854 47300 7910 47356
rect 7910 47300 7914 47356
rect 7850 47296 7914 47300
rect 12049 47356 12113 47360
rect 12049 47300 12053 47356
rect 12053 47300 12109 47356
rect 12109 47300 12113 47356
rect 12049 47296 12113 47300
rect 12129 47356 12193 47360
rect 12129 47300 12133 47356
rect 12133 47300 12189 47356
rect 12189 47300 12193 47356
rect 12129 47296 12193 47300
rect 12209 47356 12273 47360
rect 12209 47300 12213 47356
rect 12213 47300 12269 47356
rect 12269 47300 12273 47356
rect 12209 47296 12273 47300
rect 12289 47356 12353 47360
rect 12289 47300 12293 47356
rect 12293 47300 12349 47356
rect 12349 47300 12353 47356
rect 12289 47296 12353 47300
rect 16488 47356 16552 47360
rect 16488 47300 16492 47356
rect 16492 47300 16548 47356
rect 16548 47300 16552 47356
rect 16488 47296 16552 47300
rect 16568 47356 16632 47360
rect 16568 47300 16572 47356
rect 16572 47300 16628 47356
rect 16628 47300 16632 47356
rect 16568 47296 16632 47300
rect 16648 47356 16712 47360
rect 16648 47300 16652 47356
rect 16652 47300 16708 47356
rect 16708 47300 16712 47356
rect 16648 47296 16712 47300
rect 16728 47356 16792 47360
rect 16728 47300 16732 47356
rect 16732 47300 16788 47356
rect 16788 47300 16792 47356
rect 16728 47296 16792 47300
rect 5390 46812 5454 46816
rect 5390 46756 5394 46812
rect 5394 46756 5450 46812
rect 5450 46756 5454 46812
rect 5390 46752 5454 46756
rect 5470 46812 5534 46816
rect 5470 46756 5474 46812
rect 5474 46756 5530 46812
rect 5530 46756 5534 46812
rect 5470 46752 5534 46756
rect 5550 46812 5614 46816
rect 5550 46756 5554 46812
rect 5554 46756 5610 46812
rect 5610 46756 5614 46812
rect 5550 46752 5614 46756
rect 5630 46812 5694 46816
rect 5630 46756 5634 46812
rect 5634 46756 5690 46812
rect 5690 46756 5694 46812
rect 5630 46752 5694 46756
rect 9829 46812 9893 46816
rect 9829 46756 9833 46812
rect 9833 46756 9889 46812
rect 9889 46756 9893 46812
rect 9829 46752 9893 46756
rect 9909 46812 9973 46816
rect 9909 46756 9913 46812
rect 9913 46756 9969 46812
rect 9969 46756 9973 46812
rect 9909 46752 9973 46756
rect 9989 46812 10053 46816
rect 9989 46756 9993 46812
rect 9993 46756 10049 46812
rect 10049 46756 10053 46812
rect 9989 46752 10053 46756
rect 10069 46812 10133 46816
rect 10069 46756 10073 46812
rect 10073 46756 10129 46812
rect 10129 46756 10133 46812
rect 10069 46752 10133 46756
rect 14268 46812 14332 46816
rect 14268 46756 14272 46812
rect 14272 46756 14328 46812
rect 14328 46756 14332 46812
rect 14268 46752 14332 46756
rect 14348 46812 14412 46816
rect 14348 46756 14352 46812
rect 14352 46756 14408 46812
rect 14408 46756 14412 46812
rect 14348 46752 14412 46756
rect 14428 46812 14492 46816
rect 14428 46756 14432 46812
rect 14432 46756 14488 46812
rect 14488 46756 14492 46812
rect 14428 46752 14492 46756
rect 14508 46812 14572 46816
rect 14508 46756 14512 46812
rect 14512 46756 14568 46812
rect 14568 46756 14572 46812
rect 14508 46752 14572 46756
rect 18707 46812 18771 46816
rect 18707 46756 18711 46812
rect 18711 46756 18767 46812
rect 18767 46756 18771 46812
rect 18707 46752 18771 46756
rect 18787 46812 18851 46816
rect 18787 46756 18791 46812
rect 18791 46756 18847 46812
rect 18847 46756 18851 46812
rect 18787 46752 18851 46756
rect 18867 46812 18931 46816
rect 18867 46756 18871 46812
rect 18871 46756 18927 46812
rect 18927 46756 18931 46812
rect 18867 46752 18931 46756
rect 18947 46812 19011 46816
rect 18947 46756 18951 46812
rect 18951 46756 19007 46812
rect 19007 46756 19011 46812
rect 18947 46752 19011 46756
rect 3171 46268 3235 46272
rect 3171 46212 3175 46268
rect 3175 46212 3231 46268
rect 3231 46212 3235 46268
rect 3171 46208 3235 46212
rect 3251 46268 3315 46272
rect 3251 46212 3255 46268
rect 3255 46212 3311 46268
rect 3311 46212 3315 46268
rect 3251 46208 3315 46212
rect 3331 46268 3395 46272
rect 3331 46212 3335 46268
rect 3335 46212 3391 46268
rect 3391 46212 3395 46268
rect 3331 46208 3395 46212
rect 3411 46268 3475 46272
rect 3411 46212 3415 46268
rect 3415 46212 3471 46268
rect 3471 46212 3475 46268
rect 3411 46208 3475 46212
rect 7610 46268 7674 46272
rect 7610 46212 7614 46268
rect 7614 46212 7670 46268
rect 7670 46212 7674 46268
rect 7610 46208 7674 46212
rect 7690 46268 7754 46272
rect 7690 46212 7694 46268
rect 7694 46212 7750 46268
rect 7750 46212 7754 46268
rect 7690 46208 7754 46212
rect 7770 46268 7834 46272
rect 7770 46212 7774 46268
rect 7774 46212 7830 46268
rect 7830 46212 7834 46268
rect 7770 46208 7834 46212
rect 7850 46268 7914 46272
rect 7850 46212 7854 46268
rect 7854 46212 7910 46268
rect 7910 46212 7914 46268
rect 7850 46208 7914 46212
rect 12049 46268 12113 46272
rect 12049 46212 12053 46268
rect 12053 46212 12109 46268
rect 12109 46212 12113 46268
rect 12049 46208 12113 46212
rect 12129 46268 12193 46272
rect 12129 46212 12133 46268
rect 12133 46212 12189 46268
rect 12189 46212 12193 46268
rect 12129 46208 12193 46212
rect 12209 46268 12273 46272
rect 12209 46212 12213 46268
rect 12213 46212 12269 46268
rect 12269 46212 12273 46268
rect 12209 46208 12273 46212
rect 12289 46268 12353 46272
rect 12289 46212 12293 46268
rect 12293 46212 12349 46268
rect 12349 46212 12353 46268
rect 12289 46208 12353 46212
rect 16488 46268 16552 46272
rect 16488 46212 16492 46268
rect 16492 46212 16548 46268
rect 16548 46212 16552 46268
rect 16488 46208 16552 46212
rect 16568 46268 16632 46272
rect 16568 46212 16572 46268
rect 16572 46212 16628 46268
rect 16628 46212 16632 46268
rect 16568 46208 16632 46212
rect 16648 46268 16712 46272
rect 16648 46212 16652 46268
rect 16652 46212 16708 46268
rect 16708 46212 16712 46268
rect 16648 46208 16712 46212
rect 16728 46268 16792 46272
rect 16728 46212 16732 46268
rect 16732 46212 16788 46268
rect 16788 46212 16792 46268
rect 16728 46208 16792 46212
rect 5390 45724 5454 45728
rect 5390 45668 5394 45724
rect 5394 45668 5450 45724
rect 5450 45668 5454 45724
rect 5390 45664 5454 45668
rect 5470 45724 5534 45728
rect 5470 45668 5474 45724
rect 5474 45668 5530 45724
rect 5530 45668 5534 45724
rect 5470 45664 5534 45668
rect 5550 45724 5614 45728
rect 5550 45668 5554 45724
rect 5554 45668 5610 45724
rect 5610 45668 5614 45724
rect 5550 45664 5614 45668
rect 5630 45724 5694 45728
rect 5630 45668 5634 45724
rect 5634 45668 5690 45724
rect 5690 45668 5694 45724
rect 5630 45664 5694 45668
rect 9829 45724 9893 45728
rect 9829 45668 9833 45724
rect 9833 45668 9889 45724
rect 9889 45668 9893 45724
rect 9829 45664 9893 45668
rect 9909 45724 9973 45728
rect 9909 45668 9913 45724
rect 9913 45668 9969 45724
rect 9969 45668 9973 45724
rect 9909 45664 9973 45668
rect 9989 45724 10053 45728
rect 9989 45668 9993 45724
rect 9993 45668 10049 45724
rect 10049 45668 10053 45724
rect 9989 45664 10053 45668
rect 10069 45724 10133 45728
rect 10069 45668 10073 45724
rect 10073 45668 10129 45724
rect 10129 45668 10133 45724
rect 10069 45664 10133 45668
rect 14268 45724 14332 45728
rect 14268 45668 14272 45724
rect 14272 45668 14328 45724
rect 14328 45668 14332 45724
rect 14268 45664 14332 45668
rect 14348 45724 14412 45728
rect 14348 45668 14352 45724
rect 14352 45668 14408 45724
rect 14408 45668 14412 45724
rect 14348 45664 14412 45668
rect 14428 45724 14492 45728
rect 14428 45668 14432 45724
rect 14432 45668 14488 45724
rect 14488 45668 14492 45724
rect 14428 45664 14492 45668
rect 14508 45724 14572 45728
rect 14508 45668 14512 45724
rect 14512 45668 14568 45724
rect 14568 45668 14572 45724
rect 14508 45664 14572 45668
rect 18707 45724 18771 45728
rect 18707 45668 18711 45724
rect 18711 45668 18767 45724
rect 18767 45668 18771 45724
rect 18707 45664 18771 45668
rect 18787 45724 18851 45728
rect 18787 45668 18791 45724
rect 18791 45668 18847 45724
rect 18847 45668 18851 45724
rect 18787 45664 18851 45668
rect 18867 45724 18931 45728
rect 18867 45668 18871 45724
rect 18871 45668 18927 45724
rect 18927 45668 18931 45724
rect 18867 45664 18931 45668
rect 18947 45724 19011 45728
rect 18947 45668 18951 45724
rect 18951 45668 19007 45724
rect 19007 45668 19011 45724
rect 18947 45664 19011 45668
rect 3171 45180 3235 45184
rect 3171 45124 3175 45180
rect 3175 45124 3231 45180
rect 3231 45124 3235 45180
rect 3171 45120 3235 45124
rect 3251 45180 3315 45184
rect 3251 45124 3255 45180
rect 3255 45124 3311 45180
rect 3311 45124 3315 45180
rect 3251 45120 3315 45124
rect 3331 45180 3395 45184
rect 3331 45124 3335 45180
rect 3335 45124 3391 45180
rect 3391 45124 3395 45180
rect 3331 45120 3395 45124
rect 3411 45180 3475 45184
rect 3411 45124 3415 45180
rect 3415 45124 3471 45180
rect 3471 45124 3475 45180
rect 3411 45120 3475 45124
rect 7610 45180 7674 45184
rect 7610 45124 7614 45180
rect 7614 45124 7670 45180
rect 7670 45124 7674 45180
rect 7610 45120 7674 45124
rect 7690 45180 7754 45184
rect 7690 45124 7694 45180
rect 7694 45124 7750 45180
rect 7750 45124 7754 45180
rect 7690 45120 7754 45124
rect 7770 45180 7834 45184
rect 7770 45124 7774 45180
rect 7774 45124 7830 45180
rect 7830 45124 7834 45180
rect 7770 45120 7834 45124
rect 7850 45180 7914 45184
rect 7850 45124 7854 45180
rect 7854 45124 7910 45180
rect 7910 45124 7914 45180
rect 7850 45120 7914 45124
rect 12049 45180 12113 45184
rect 12049 45124 12053 45180
rect 12053 45124 12109 45180
rect 12109 45124 12113 45180
rect 12049 45120 12113 45124
rect 12129 45180 12193 45184
rect 12129 45124 12133 45180
rect 12133 45124 12189 45180
rect 12189 45124 12193 45180
rect 12129 45120 12193 45124
rect 12209 45180 12273 45184
rect 12209 45124 12213 45180
rect 12213 45124 12269 45180
rect 12269 45124 12273 45180
rect 12209 45120 12273 45124
rect 12289 45180 12353 45184
rect 12289 45124 12293 45180
rect 12293 45124 12349 45180
rect 12349 45124 12353 45180
rect 12289 45120 12353 45124
rect 16488 45180 16552 45184
rect 16488 45124 16492 45180
rect 16492 45124 16548 45180
rect 16548 45124 16552 45180
rect 16488 45120 16552 45124
rect 16568 45180 16632 45184
rect 16568 45124 16572 45180
rect 16572 45124 16628 45180
rect 16628 45124 16632 45180
rect 16568 45120 16632 45124
rect 16648 45180 16712 45184
rect 16648 45124 16652 45180
rect 16652 45124 16708 45180
rect 16708 45124 16712 45180
rect 16648 45120 16712 45124
rect 16728 45180 16792 45184
rect 16728 45124 16732 45180
rect 16732 45124 16788 45180
rect 16788 45124 16792 45180
rect 16728 45120 16792 45124
rect 5390 44636 5454 44640
rect 5390 44580 5394 44636
rect 5394 44580 5450 44636
rect 5450 44580 5454 44636
rect 5390 44576 5454 44580
rect 5470 44636 5534 44640
rect 5470 44580 5474 44636
rect 5474 44580 5530 44636
rect 5530 44580 5534 44636
rect 5470 44576 5534 44580
rect 5550 44636 5614 44640
rect 5550 44580 5554 44636
rect 5554 44580 5610 44636
rect 5610 44580 5614 44636
rect 5550 44576 5614 44580
rect 5630 44636 5694 44640
rect 5630 44580 5634 44636
rect 5634 44580 5690 44636
rect 5690 44580 5694 44636
rect 5630 44576 5694 44580
rect 9829 44636 9893 44640
rect 9829 44580 9833 44636
rect 9833 44580 9889 44636
rect 9889 44580 9893 44636
rect 9829 44576 9893 44580
rect 9909 44636 9973 44640
rect 9909 44580 9913 44636
rect 9913 44580 9969 44636
rect 9969 44580 9973 44636
rect 9909 44576 9973 44580
rect 9989 44636 10053 44640
rect 9989 44580 9993 44636
rect 9993 44580 10049 44636
rect 10049 44580 10053 44636
rect 9989 44576 10053 44580
rect 10069 44636 10133 44640
rect 10069 44580 10073 44636
rect 10073 44580 10129 44636
rect 10129 44580 10133 44636
rect 10069 44576 10133 44580
rect 14268 44636 14332 44640
rect 14268 44580 14272 44636
rect 14272 44580 14328 44636
rect 14328 44580 14332 44636
rect 14268 44576 14332 44580
rect 14348 44636 14412 44640
rect 14348 44580 14352 44636
rect 14352 44580 14408 44636
rect 14408 44580 14412 44636
rect 14348 44576 14412 44580
rect 14428 44636 14492 44640
rect 14428 44580 14432 44636
rect 14432 44580 14488 44636
rect 14488 44580 14492 44636
rect 14428 44576 14492 44580
rect 14508 44636 14572 44640
rect 14508 44580 14512 44636
rect 14512 44580 14568 44636
rect 14568 44580 14572 44636
rect 14508 44576 14572 44580
rect 18707 44636 18771 44640
rect 18707 44580 18711 44636
rect 18711 44580 18767 44636
rect 18767 44580 18771 44636
rect 18707 44576 18771 44580
rect 18787 44636 18851 44640
rect 18787 44580 18791 44636
rect 18791 44580 18847 44636
rect 18847 44580 18851 44636
rect 18787 44576 18851 44580
rect 18867 44636 18931 44640
rect 18867 44580 18871 44636
rect 18871 44580 18927 44636
rect 18927 44580 18931 44636
rect 18867 44576 18931 44580
rect 18947 44636 19011 44640
rect 18947 44580 18951 44636
rect 18951 44580 19007 44636
rect 19007 44580 19011 44636
rect 18947 44576 19011 44580
rect 3171 44092 3235 44096
rect 3171 44036 3175 44092
rect 3175 44036 3231 44092
rect 3231 44036 3235 44092
rect 3171 44032 3235 44036
rect 3251 44092 3315 44096
rect 3251 44036 3255 44092
rect 3255 44036 3311 44092
rect 3311 44036 3315 44092
rect 3251 44032 3315 44036
rect 3331 44092 3395 44096
rect 3331 44036 3335 44092
rect 3335 44036 3391 44092
rect 3391 44036 3395 44092
rect 3331 44032 3395 44036
rect 3411 44092 3475 44096
rect 3411 44036 3415 44092
rect 3415 44036 3471 44092
rect 3471 44036 3475 44092
rect 3411 44032 3475 44036
rect 7610 44092 7674 44096
rect 7610 44036 7614 44092
rect 7614 44036 7670 44092
rect 7670 44036 7674 44092
rect 7610 44032 7674 44036
rect 7690 44092 7754 44096
rect 7690 44036 7694 44092
rect 7694 44036 7750 44092
rect 7750 44036 7754 44092
rect 7690 44032 7754 44036
rect 7770 44092 7834 44096
rect 7770 44036 7774 44092
rect 7774 44036 7830 44092
rect 7830 44036 7834 44092
rect 7770 44032 7834 44036
rect 7850 44092 7914 44096
rect 7850 44036 7854 44092
rect 7854 44036 7910 44092
rect 7910 44036 7914 44092
rect 7850 44032 7914 44036
rect 12049 44092 12113 44096
rect 12049 44036 12053 44092
rect 12053 44036 12109 44092
rect 12109 44036 12113 44092
rect 12049 44032 12113 44036
rect 12129 44092 12193 44096
rect 12129 44036 12133 44092
rect 12133 44036 12189 44092
rect 12189 44036 12193 44092
rect 12129 44032 12193 44036
rect 12209 44092 12273 44096
rect 12209 44036 12213 44092
rect 12213 44036 12269 44092
rect 12269 44036 12273 44092
rect 12209 44032 12273 44036
rect 12289 44092 12353 44096
rect 12289 44036 12293 44092
rect 12293 44036 12349 44092
rect 12349 44036 12353 44092
rect 12289 44032 12353 44036
rect 16488 44092 16552 44096
rect 16488 44036 16492 44092
rect 16492 44036 16548 44092
rect 16548 44036 16552 44092
rect 16488 44032 16552 44036
rect 16568 44092 16632 44096
rect 16568 44036 16572 44092
rect 16572 44036 16628 44092
rect 16628 44036 16632 44092
rect 16568 44032 16632 44036
rect 16648 44092 16712 44096
rect 16648 44036 16652 44092
rect 16652 44036 16708 44092
rect 16708 44036 16712 44092
rect 16648 44032 16712 44036
rect 16728 44092 16792 44096
rect 16728 44036 16732 44092
rect 16732 44036 16788 44092
rect 16788 44036 16792 44092
rect 16728 44032 16792 44036
rect 5390 43548 5454 43552
rect 5390 43492 5394 43548
rect 5394 43492 5450 43548
rect 5450 43492 5454 43548
rect 5390 43488 5454 43492
rect 5470 43548 5534 43552
rect 5470 43492 5474 43548
rect 5474 43492 5530 43548
rect 5530 43492 5534 43548
rect 5470 43488 5534 43492
rect 5550 43548 5614 43552
rect 5550 43492 5554 43548
rect 5554 43492 5610 43548
rect 5610 43492 5614 43548
rect 5550 43488 5614 43492
rect 5630 43548 5694 43552
rect 5630 43492 5634 43548
rect 5634 43492 5690 43548
rect 5690 43492 5694 43548
rect 5630 43488 5694 43492
rect 9829 43548 9893 43552
rect 9829 43492 9833 43548
rect 9833 43492 9889 43548
rect 9889 43492 9893 43548
rect 9829 43488 9893 43492
rect 9909 43548 9973 43552
rect 9909 43492 9913 43548
rect 9913 43492 9969 43548
rect 9969 43492 9973 43548
rect 9909 43488 9973 43492
rect 9989 43548 10053 43552
rect 9989 43492 9993 43548
rect 9993 43492 10049 43548
rect 10049 43492 10053 43548
rect 9989 43488 10053 43492
rect 10069 43548 10133 43552
rect 10069 43492 10073 43548
rect 10073 43492 10129 43548
rect 10129 43492 10133 43548
rect 10069 43488 10133 43492
rect 14268 43548 14332 43552
rect 14268 43492 14272 43548
rect 14272 43492 14328 43548
rect 14328 43492 14332 43548
rect 14268 43488 14332 43492
rect 14348 43548 14412 43552
rect 14348 43492 14352 43548
rect 14352 43492 14408 43548
rect 14408 43492 14412 43548
rect 14348 43488 14412 43492
rect 14428 43548 14492 43552
rect 14428 43492 14432 43548
rect 14432 43492 14488 43548
rect 14488 43492 14492 43548
rect 14428 43488 14492 43492
rect 14508 43548 14572 43552
rect 14508 43492 14512 43548
rect 14512 43492 14568 43548
rect 14568 43492 14572 43548
rect 14508 43488 14572 43492
rect 18707 43548 18771 43552
rect 18707 43492 18711 43548
rect 18711 43492 18767 43548
rect 18767 43492 18771 43548
rect 18707 43488 18771 43492
rect 18787 43548 18851 43552
rect 18787 43492 18791 43548
rect 18791 43492 18847 43548
rect 18847 43492 18851 43548
rect 18787 43488 18851 43492
rect 18867 43548 18931 43552
rect 18867 43492 18871 43548
rect 18871 43492 18927 43548
rect 18927 43492 18931 43548
rect 18867 43488 18931 43492
rect 18947 43548 19011 43552
rect 18947 43492 18951 43548
rect 18951 43492 19007 43548
rect 19007 43492 19011 43548
rect 18947 43488 19011 43492
rect 3171 43004 3235 43008
rect 3171 42948 3175 43004
rect 3175 42948 3231 43004
rect 3231 42948 3235 43004
rect 3171 42944 3235 42948
rect 3251 43004 3315 43008
rect 3251 42948 3255 43004
rect 3255 42948 3311 43004
rect 3311 42948 3315 43004
rect 3251 42944 3315 42948
rect 3331 43004 3395 43008
rect 3331 42948 3335 43004
rect 3335 42948 3391 43004
rect 3391 42948 3395 43004
rect 3331 42944 3395 42948
rect 3411 43004 3475 43008
rect 3411 42948 3415 43004
rect 3415 42948 3471 43004
rect 3471 42948 3475 43004
rect 3411 42944 3475 42948
rect 7610 43004 7674 43008
rect 7610 42948 7614 43004
rect 7614 42948 7670 43004
rect 7670 42948 7674 43004
rect 7610 42944 7674 42948
rect 7690 43004 7754 43008
rect 7690 42948 7694 43004
rect 7694 42948 7750 43004
rect 7750 42948 7754 43004
rect 7690 42944 7754 42948
rect 7770 43004 7834 43008
rect 7770 42948 7774 43004
rect 7774 42948 7830 43004
rect 7830 42948 7834 43004
rect 7770 42944 7834 42948
rect 7850 43004 7914 43008
rect 7850 42948 7854 43004
rect 7854 42948 7910 43004
rect 7910 42948 7914 43004
rect 7850 42944 7914 42948
rect 12049 43004 12113 43008
rect 12049 42948 12053 43004
rect 12053 42948 12109 43004
rect 12109 42948 12113 43004
rect 12049 42944 12113 42948
rect 12129 43004 12193 43008
rect 12129 42948 12133 43004
rect 12133 42948 12189 43004
rect 12189 42948 12193 43004
rect 12129 42944 12193 42948
rect 12209 43004 12273 43008
rect 12209 42948 12213 43004
rect 12213 42948 12269 43004
rect 12269 42948 12273 43004
rect 12209 42944 12273 42948
rect 12289 43004 12353 43008
rect 12289 42948 12293 43004
rect 12293 42948 12349 43004
rect 12349 42948 12353 43004
rect 12289 42944 12353 42948
rect 16488 43004 16552 43008
rect 16488 42948 16492 43004
rect 16492 42948 16548 43004
rect 16548 42948 16552 43004
rect 16488 42944 16552 42948
rect 16568 43004 16632 43008
rect 16568 42948 16572 43004
rect 16572 42948 16628 43004
rect 16628 42948 16632 43004
rect 16568 42944 16632 42948
rect 16648 43004 16712 43008
rect 16648 42948 16652 43004
rect 16652 42948 16708 43004
rect 16708 42948 16712 43004
rect 16648 42944 16712 42948
rect 16728 43004 16792 43008
rect 16728 42948 16732 43004
rect 16732 42948 16788 43004
rect 16788 42948 16792 43004
rect 16728 42944 16792 42948
rect 5390 42460 5454 42464
rect 5390 42404 5394 42460
rect 5394 42404 5450 42460
rect 5450 42404 5454 42460
rect 5390 42400 5454 42404
rect 5470 42460 5534 42464
rect 5470 42404 5474 42460
rect 5474 42404 5530 42460
rect 5530 42404 5534 42460
rect 5470 42400 5534 42404
rect 5550 42460 5614 42464
rect 5550 42404 5554 42460
rect 5554 42404 5610 42460
rect 5610 42404 5614 42460
rect 5550 42400 5614 42404
rect 5630 42460 5694 42464
rect 5630 42404 5634 42460
rect 5634 42404 5690 42460
rect 5690 42404 5694 42460
rect 5630 42400 5694 42404
rect 9829 42460 9893 42464
rect 9829 42404 9833 42460
rect 9833 42404 9889 42460
rect 9889 42404 9893 42460
rect 9829 42400 9893 42404
rect 9909 42460 9973 42464
rect 9909 42404 9913 42460
rect 9913 42404 9969 42460
rect 9969 42404 9973 42460
rect 9909 42400 9973 42404
rect 9989 42460 10053 42464
rect 9989 42404 9993 42460
rect 9993 42404 10049 42460
rect 10049 42404 10053 42460
rect 9989 42400 10053 42404
rect 10069 42460 10133 42464
rect 10069 42404 10073 42460
rect 10073 42404 10129 42460
rect 10129 42404 10133 42460
rect 10069 42400 10133 42404
rect 14268 42460 14332 42464
rect 14268 42404 14272 42460
rect 14272 42404 14328 42460
rect 14328 42404 14332 42460
rect 14268 42400 14332 42404
rect 14348 42460 14412 42464
rect 14348 42404 14352 42460
rect 14352 42404 14408 42460
rect 14408 42404 14412 42460
rect 14348 42400 14412 42404
rect 14428 42460 14492 42464
rect 14428 42404 14432 42460
rect 14432 42404 14488 42460
rect 14488 42404 14492 42460
rect 14428 42400 14492 42404
rect 14508 42460 14572 42464
rect 14508 42404 14512 42460
rect 14512 42404 14568 42460
rect 14568 42404 14572 42460
rect 14508 42400 14572 42404
rect 18707 42460 18771 42464
rect 18707 42404 18711 42460
rect 18711 42404 18767 42460
rect 18767 42404 18771 42460
rect 18707 42400 18771 42404
rect 18787 42460 18851 42464
rect 18787 42404 18791 42460
rect 18791 42404 18847 42460
rect 18847 42404 18851 42460
rect 18787 42400 18851 42404
rect 18867 42460 18931 42464
rect 18867 42404 18871 42460
rect 18871 42404 18927 42460
rect 18927 42404 18931 42460
rect 18867 42400 18931 42404
rect 18947 42460 19011 42464
rect 18947 42404 18951 42460
rect 18951 42404 19007 42460
rect 19007 42404 19011 42460
rect 18947 42400 19011 42404
rect 3171 41916 3235 41920
rect 3171 41860 3175 41916
rect 3175 41860 3231 41916
rect 3231 41860 3235 41916
rect 3171 41856 3235 41860
rect 3251 41916 3315 41920
rect 3251 41860 3255 41916
rect 3255 41860 3311 41916
rect 3311 41860 3315 41916
rect 3251 41856 3315 41860
rect 3331 41916 3395 41920
rect 3331 41860 3335 41916
rect 3335 41860 3391 41916
rect 3391 41860 3395 41916
rect 3331 41856 3395 41860
rect 3411 41916 3475 41920
rect 3411 41860 3415 41916
rect 3415 41860 3471 41916
rect 3471 41860 3475 41916
rect 3411 41856 3475 41860
rect 7610 41916 7674 41920
rect 7610 41860 7614 41916
rect 7614 41860 7670 41916
rect 7670 41860 7674 41916
rect 7610 41856 7674 41860
rect 7690 41916 7754 41920
rect 7690 41860 7694 41916
rect 7694 41860 7750 41916
rect 7750 41860 7754 41916
rect 7690 41856 7754 41860
rect 7770 41916 7834 41920
rect 7770 41860 7774 41916
rect 7774 41860 7830 41916
rect 7830 41860 7834 41916
rect 7770 41856 7834 41860
rect 7850 41916 7914 41920
rect 7850 41860 7854 41916
rect 7854 41860 7910 41916
rect 7910 41860 7914 41916
rect 7850 41856 7914 41860
rect 12049 41916 12113 41920
rect 12049 41860 12053 41916
rect 12053 41860 12109 41916
rect 12109 41860 12113 41916
rect 12049 41856 12113 41860
rect 12129 41916 12193 41920
rect 12129 41860 12133 41916
rect 12133 41860 12189 41916
rect 12189 41860 12193 41916
rect 12129 41856 12193 41860
rect 12209 41916 12273 41920
rect 12209 41860 12213 41916
rect 12213 41860 12269 41916
rect 12269 41860 12273 41916
rect 12209 41856 12273 41860
rect 12289 41916 12353 41920
rect 12289 41860 12293 41916
rect 12293 41860 12349 41916
rect 12349 41860 12353 41916
rect 12289 41856 12353 41860
rect 16488 41916 16552 41920
rect 16488 41860 16492 41916
rect 16492 41860 16548 41916
rect 16548 41860 16552 41916
rect 16488 41856 16552 41860
rect 16568 41916 16632 41920
rect 16568 41860 16572 41916
rect 16572 41860 16628 41916
rect 16628 41860 16632 41916
rect 16568 41856 16632 41860
rect 16648 41916 16712 41920
rect 16648 41860 16652 41916
rect 16652 41860 16708 41916
rect 16708 41860 16712 41916
rect 16648 41856 16712 41860
rect 16728 41916 16792 41920
rect 16728 41860 16732 41916
rect 16732 41860 16788 41916
rect 16788 41860 16792 41916
rect 16728 41856 16792 41860
rect 5390 41372 5454 41376
rect 5390 41316 5394 41372
rect 5394 41316 5450 41372
rect 5450 41316 5454 41372
rect 5390 41312 5454 41316
rect 5470 41372 5534 41376
rect 5470 41316 5474 41372
rect 5474 41316 5530 41372
rect 5530 41316 5534 41372
rect 5470 41312 5534 41316
rect 5550 41372 5614 41376
rect 5550 41316 5554 41372
rect 5554 41316 5610 41372
rect 5610 41316 5614 41372
rect 5550 41312 5614 41316
rect 5630 41372 5694 41376
rect 5630 41316 5634 41372
rect 5634 41316 5690 41372
rect 5690 41316 5694 41372
rect 5630 41312 5694 41316
rect 9829 41372 9893 41376
rect 9829 41316 9833 41372
rect 9833 41316 9889 41372
rect 9889 41316 9893 41372
rect 9829 41312 9893 41316
rect 9909 41372 9973 41376
rect 9909 41316 9913 41372
rect 9913 41316 9969 41372
rect 9969 41316 9973 41372
rect 9909 41312 9973 41316
rect 9989 41372 10053 41376
rect 9989 41316 9993 41372
rect 9993 41316 10049 41372
rect 10049 41316 10053 41372
rect 9989 41312 10053 41316
rect 10069 41372 10133 41376
rect 10069 41316 10073 41372
rect 10073 41316 10129 41372
rect 10129 41316 10133 41372
rect 10069 41312 10133 41316
rect 14268 41372 14332 41376
rect 14268 41316 14272 41372
rect 14272 41316 14328 41372
rect 14328 41316 14332 41372
rect 14268 41312 14332 41316
rect 14348 41372 14412 41376
rect 14348 41316 14352 41372
rect 14352 41316 14408 41372
rect 14408 41316 14412 41372
rect 14348 41312 14412 41316
rect 14428 41372 14492 41376
rect 14428 41316 14432 41372
rect 14432 41316 14488 41372
rect 14488 41316 14492 41372
rect 14428 41312 14492 41316
rect 14508 41372 14572 41376
rect 14508 41316 14512 41372
rect 14512 41316 14568 41372
rect 14568 41316 14572 41372
rect 14508 41312 14572 41316
rect 18707 41372 18771 41376
rect 18707 41316 18711 41372
rect 18711 41316 18767 41372
rect 18767 41316 18771 41372
rect 18707 41312 18771 41316
rect 18787 41372 18851 41376
rect 18787 41316 18791 41372
rect 18791 41316 18847 41372
rect 18847 41316 18851 41372
rect 18787 41312 18851 41316
rect 18867 41372 18931 41376
rect 18867 41316 18871 41372
rect 18871 41316 18927 41372
rect 18927 41316 18931 41372
rect 18867 41312 18931 41316
rect 18947 41372 19011 41376
rect 18947 41316 18951 41372
rect 18951 41316 19007 41372
rect 19007 41316 19011 41372
rect 18947 41312 19011 41316
rect 3171 40828 3235 40832
rect 3171 40772 3175 40828
rect 3175 40772 3231 40828
rect 3231 40772 3235 40828
rect 3171 40768 3235 40772
rect 3251 40828 3315 40832
rect 3251 40772 3255 40828
rect 3255 40772 3311 40828
rect 3311 40772 3315 40828
rect 3251 40768 3315 40772
rect 3331 40828 3395 40832
rect 3331 40772 3335 40828
rect 3335 40772 3391 40828
rect 3391 40772 3395 40828
rect 3331 40768 3395 40772
rect 3411 40828 3475 40832
rect 3411 40772 3415 40828
rect 3415 40772 3471 40828
rect 3471 40772 3475 40828
rect 3411 40768 3475 40772
rect 7610 40828 7674 40832
rect 7610 40772 7614 40828
rect 7614 40772 7670 40828
rect 7670 40772 7674 40828
rect 7610 40768 7674 40772
rect 7690 40828 7754 40832
rect 7690 40772 7694 40828
rect 7694 40772 7750 40828
rect 7750 40772 7754 40828
rect 7690 40768 7754 40772
rect 7770 40828 7834 40832
rect 7770 40772 7774 40828
rect 7774 40772 7830 40828
rect 7830 40772 7834 40828
rect 7770 40768 7834 40772
rect 7850 40828 7914 40832
rect 7850 40772 7854 40828
rect 7854 40772 7910 40828
rect 7910 40772 7914 40828
rect 7850 40768 7914 40772
rect 12049 40828 12113 40832
rect 12049 40772 12053 40828
rect 12053 40772 12109 40828
rect 12109 40772 12113 40828
rect 12049 40768 12113 40772
rect 12129 40828 12193 40832
rect 12129 40772 12133 40828
rect 12133 40772 12189 40828
rect 12189 40772 12193 40828
rect 12129 40768 12193 40772
rect 12209 40828 12273 40832
rect 12209 40772 12213 40828
rect 12213 40772 12269 40828
rect 12269 40772 12273 40828
rect 12209 40768 12273 40772
rect 12289 40828 12353 40832
rect 12289 40772 12293 40828
rect 12293 40772 12349 40828
rect 12349 40772 12353 40828
rect 12289 40768 12353 40772
rect 16488 40828 16552 40832
rect 16488 40772 16492 40828
rect 16492 40772 16548 40828
rect 16548 40772 16552 40828
rect 16488 40768 16552 40772
rect 16568 40828 16632 40832
rect 16568 40772 16572 40828
rect 16572 40772 16628 40828
rect 16628 40772 16632 40828
rect 16568 40768 16632 40772
rect 16648 40828 16712 40832
rect 16648 40772 16652 40828
rect 16652 40772 16708 40828
rect 16708 40772 16712 40828
rect 16648 40768 16712 40772
rect 16728 40828 16792 40832
rect 16728 40772 16732 40828
rect 16732 40772 16788 40828
rect 16788 40772 16792 40828
rect 16728 40768 16792 40772
rect 5390 40284 5454 40288
rect 5390 40228 5394 40284
rect 5394 40228 5450 40284
rect 5450 40228 5454 40284
rect 5390 40224 5454 40228
rect 5470 40284 5534 40288
rect 5470 40228 5474 40284
rect 5474 40228 5530 40284
rect 5530 40228 5534 40284
rect 5470 40224 5534 40228
rect 5550 40284 5614 40288
rect 5550 40228 5554 40284
rect 5554 40228 5610 40284
rect 5610 40228 5614 40284
rect 5550 40224 5614 40228
rect 5630 40284 5694 40288
rect 5630 40228 5634 40284
rect 5634 40228 5690 40284
rect 5690 40228 5694 40284
rect 5630 40224 5694 40228
rect 9829 40284 9893 40288
rect 9829 40228 9833 40284
rect 9833 40228 9889 40284
rect 9889 40228 9893 40284
rect 9829 40224 9893 40228
rect 9909 40284 9973 40288
rect 9909 40228 9913 40284
rect 9913 40228 9969 40284
rect 9969 40228 9973 40284
rect 9909 40224 9973 40228
rect 9989 40284 10053 40288
rect 9989 40228 9993 40284
rect 9993 40228 10049 40284
rect 10049 40228 10053 40284
rect 9989 40224 10053 40228
rect 10069 40284 10133 40288
rect 10069 40228 10073 40284
rect 10073 40228 10129 40284
rect 10129 40228 10133 40284
rect 10069 40224 10133 40228
rect 14268 40284 14332 40288
rect 14268 40228 14272 40284
rect 14272 40228 14328 40284
rect 14328 40228 14332 40284
rect 14268 40224 14332 40228
rect 14348 40284 14412 40288
rect 14348 40228 14352 40284
rect 14352 40228 14408 40284
rect 14408 40228 14412 40284
rect 14348 40224 14412 40228
rect 14428 40284 14492 40288
rect 14428 40228 14432 40284
rect 14432 40228 14488 40284
rect 14488 40228 14492 40284
rect 14428 40224 14492 40228
rect 14508 40284 14572 40288
rect 14508 40228 14512 40284
rect 14512 40228 14568 40284
rect 14568 40228 14572 40284
rect 14508 40224 14572 40228
rect 18707 40284 18771 40288
rect 18707 40228 18711 40284
rect 18711 40228 18767 40284
rect 18767 40228 18771 40284
rect 18707 40224 18771 40228
rect 18787 40284 18851 40288
rect 18787 40228 18791 40284
rect 18791 40228 18847 40284
rect 18847 40228 18851 40284
rect 18787 40224 18851 40228
rect 18867 40284 18931 40288
rect 18867 40228 18871 40284
rect 18871 40228 18927 40284
rect 18927 40228 18931 40284
rect 18867 40224 18931 40228
rect 18947 40284 19011 40288
rect 18947 40228 18951 40284
rect 18951 40228 19007 40284
rect 19007 40228 19011 40284
rect 18947 40224 19011 40228
rect 3171 39740 3235 39744
rect 3171 39684 3175 39740
rect 3175 39684 3231 39740
rect 3231 39684 3235 39740
rect 3171 39680 3235 39684
rect 3251 39740 3315 39744
rect 3251 39684 3255 39740
rect 3255 39684 3311 39740
rect 3311 39684 3315 39740
rect 3251 39680 3315 39684
rect 3331 39740 3395 39744
rect 3331 39684 3335 39740
rect 3335 39684 3391 39740
rect 3391 39684 3395 39740
rect 3331 39680 3395 39684
rect 3411 39740 3475 39744
rect 3411 39684 3415 39740
rect 3415 39684 3471 39740
rect 3471 39684 3475 39740
rect 3411 39680 3475 39684
rect 7610 39740 7674 39744
rect 7610 39684 7614 39740
rect 7614 39684 7670 39740
rect 7670 39684 7674 39740
rect 7610 39680 7674 39684
rect 7690 39740 7754 39744
rect 7690 39684 7694 39740
rect 7694 39684 7750 39740
rect 7750 39684 7754 39740
rect 7690 39680 7754 39684
rect 7770 39740 7834 39744
rect 7770 39684 7774 39740
rect 7774 39684 7830 39740
rect 7830 39684 7834 39740
rect 7770 39680 7834 39684
rect 7850 39740 7914 39744
rect 7850 39684 7854 39740
rect 7854 39684 7910 39740
rect 7910 39684 7914 39740
rect 7850 39680 7914 39684
rect 12049 39740 12113 39744
rect 12049 39684 12053 39740
rect 12053 39684 12109 39740
rect 12109 39684 12113 39740
rect 12049 39680 12113 39684
rect 12129 39740 12193 39744
rect 12129 39684 12133 39740
rect 12133 39684 12189 39740
rect 12189 39684 12193 39740
rect 12129 39680 12193 39684
rect 12209 39740 12273 39744
rect 12209 39684 12213 39740
rect 12213 39684 12269 39740
rect 12269 39684 12273 39740
rect 12209 39680 12273 39684
rect 12289 39740 12353 39744
rect 12289 39684 12293 39740
rect 12293 39684 12349 39740
rect 12349 39684 12353 39740
rect 12289 39680 12353 39684
rect 16488 39740 16552 39744
rect 16488 39684 16492 39740
rect 16492 39684 16548 39740
rect 16548 39684 16552 39740
rect 16488 39680 16552 39684
rect 16568 39740 16632 39744
rect 16568 39684 16572 39740
rect 16572 39684 16628 39740
rect 16628 39684 16632 39740
rect 16568 39680 16632 39684
rect 16648 39740 16712 39744
rect 16648 39684 16652 39740
rect 16652 39684 16708 39740
rect 16708 39684 16712 39740
rect 16648 39680 16712 39684
rect 16728 39740 16792 39744
rect 16728 39684 16732 39740
rect 16732 39684 16788 39740
rect 16788 39684 16792 39740
rect 16728 39680 16792 39684
rect 5390 39196 5454 39200
rect 5390 39140 5394 39196
rect 5394 39140 5450 39196
rect 5450 39140 5454 39196
rect 5390 39136 5454 39140
rect 5470 39196 5534 39200
rect 5470 39140 5474 39196
rect 5474 39140 5530 39196
rect 5530 39140 5534 39196
rect 5470 39136 5534 39140
rect 5550 39196 5614 39200
rect 5550 39140 5554 39196
rect 5554 39140 5610 39196
rect 5610 39140 5614 39196
rect 5550 39136 5614 39140
rect 5630 39196 5694 39200
rect 5630 39140 5634 39196
rect 5634 39140 5690 39196
rect 5690 39140 5694 39196
rect 5630 39136 5694 39140
rect 9829 39196 9893 39200
rect 9829 39140 9833 39196
rect 9833 39140 9889 39196
rect 9889 39140 9893 39196
rect 9829 39136 9893 39140
rect 9909 39196 9973 39200
rect 9909 39140 9913 39196
rect 9913 39140 9969 39196
rect 9969 39140 9973 39196
rect 9909 39136 9973 39140
rect 9989 39196 10053 39200
rect 9989 39140 9993 39196
rect 9993 39140 10049 39196
rect 10049 39140 10053 39196
rect 9989 39136 10053 39140
rect 10069 39196 10133 39200
rect 10069 39140 10073 39196
rect 10073 39140 10129 39196
rect 10129 39140 10133 39196
rect 10069 39136 10133 39140
rect 14268 39196 14332 39200
rect 14268 39140 14272 39196
rect 14272 39140 14328 39196
rect 14328 39140 14332 39196
rect 14268 39136 14332 39140
rect 14348 39196 14412 39200
rect 14348 39140 14352 39196
rect 14352 39140 14408 39196
rect 14408 39140 14412 39196
rect 14348 39136 14412 39140
rect 14428 39196 14492 39200
rect 14428 39140 14432 39196
rect 14432 39140 14488 39196
rect 14488 39140 14492 39196
rect 14428 39136 14492 39140
rect 14508 39196 14572 39200
rect 14508 39140 14512 39196
rect 14512 39140 14568 39196
rect 14568 39140 14572 39196
rect 14508 39136 14572 39140
rect 18707 39196 18771 39200
rect 18707 39140 18711 39196
rect 18711 39140 18767 39196
rect 18767 39140 18771 39196
rect 18707 39136 18771 39140
rect 18787 39196 18851 39200
rect 18787 39140 18791 39196
rect 18791 39140 18847 39196
rect 18847 39140 18851 39196
rect 18787 39136 18851 39140
rect 18867 39196 18931 39200
rect 18867 39140 18871 39196
rect 18871 39140 18927 39196
rect 18927 39140 18931 39196
rect 18867 39136 18931 39140
rect 18947 39196 19011 39200
rect 18947 39140 18951 39196
rect 18951 39140 19007 39196
rect 19007 39140 19011 39196
rect 18947 39136 19011 39140
rect 3171 38652 3235 38656
rect 3171 38596 3175 38652
rect 3175 38596 3231 38652
rect 3231 38596 3235 38652
rect 3171 38592 3235 38596
rect 3251 38652 3315 38656
rect 3251 38596 3255 38652
rect 3255 38596 3311 38652
rect 3311 38596 3315 38652
rect 3251 38592 3315 38596
rect 3331 38652 3395 38656
rect 3331 38596 3335 38652
rect 3335 38596 3391 38652
rect 3391 38596 3395 38652
rect 3331 38592 3395 38596
rect 3411 38652 3475 38656
rect 3411 38596 3415 38652
rect 3415 38596 3471 38652
rect 3471 38596 3475 38652
rect 3411 38592 3475 38596
rect 7610 38652 7674 38656
rect 7610 38596 7614 38652
rect 7614 38596 7670 38652
rect 7670 38596 7674 38652
rect 7610 38592 7674 38596
rect 7690 38652 7754 38656
rect 7690 38596 7694 38652
rect 7694 38596 7750 38652
rect 7750 38596 7754 38652
rect 7690 38592 7754 38596
rect 7770 38652 7834 38656
rect 7770 38596 7774 38652
rect 7774 38596 7830 38652
rect 7830 38596 7834 38652
rect 7770 38592 7834 38596
rect 7850 38652 7914 38656
rect 7850 38596 7854 38652
rect 7854 38596 7910 38652
rect 7910 38596 7914 38652
rect 7850 38592 7914 38596
rect 12049 38652 12113 38656
rect 12049 38596 12053 38652
rect 12053 38596 12109 38652
rect 12109 38596 12113 38652
rect 12049 38592 12113 38596
rect 12129 38652 12193 38656
rect 12129 38596 12133 38652
rect 12133 38596 12189 38652
rect 12189 38596 12193 38652
rect 12129 38592 12193 38596
rect 12209 38652 12273 38656
rect 12209 38596 12213 38652
rect 12213 38596 12269 38652
rect 12269 38596 12273 38652
rect 12209 38592 12273 38596
rect 12289 38652 12353 38656
rect 12289 38596 12293 38652
rect 12293 38596 12349 38652
rect 12349 38596 12353 38652
rect 12289 38592 12353 38596
rect 16488 38652 16552 38656
rect 16488 38596 16492 38652
rect 16492 38596 16548 38652
rect 16548 38596 16552 38652
rect 16488 38592 16552 38596
rect 16568 38652 16632 38656
rect 16568 38596 16572 38652
rect 16572 38596 16628 38652
rect 16628 38596 16632 38652
rect 16568 38592 16632 38596
rect 16648 38652 16712 38656
rect 16648 38596 16652 38652
rect 16652 38596 16708 38652
rect 16708 38596 16712 38652
rect 16648 38592 16712 38596
rect 16728 38652 16792 38656
rect 16728 38596 16732 38652
rect 16732 38596 16788 38652
rect 16788 38596 16792 38652
rect 16728 38592 16792 38596
rect 5390 38108 5454 38112
rect 5390 38052 5394 38108
rect 5394 38052 5450 38108
rect 5450 38052 5454 38108
rect 5390 38048 5454 38052
rect 5470 38108 5534 38112
rect 5470 38052 5474 38108
rect 5474 38052 5530 38108
rect 5530 38052 5534 38108
rect 5470 38048 5534 38052
rect 5550 38108 5614 38112
rect 5550 38052 5554 38108
rect 5554 38052 5610 38108
rect 5610 38052 5614 38108
rect 5550 38048 5614 38052
rect 5630 38108 5694 38112
rect 5630 38052 5634 38108
rect 5634 38052 5690 38108
rect 5690 38052 5694 38108
rect 5630 38048 5694 38052
rect 9829 38108 9893 38112
rect 9829 38052 9833 38108
rect 9833 38052 9889 38108
rect 9889 38052 9893 38108
rect 9829 38048 9893 38052
rect 9909 38108 9973 38112
rect 9909 38052 9913 38108
rect 9913 38052 9969 38108
rect 9969 38052 9973 38108
rect 9909 38048 9973 38052
rect 9989 38108 10053 38112
rect 9989 38052 9993 38108
rect 9993 38052 10049 38108
rect 10049 38052 10053 38108
rect 9989 38048 10053 38052
rect 10069 38108 10133 38112
rect 10069 38052 10073 38108
rect 10073 38052 10129 38108
rect 10129 38052 10133 38108
rect 10069 38048 10133 38052
rect 14268 38108 14332 38112
rect 14268 38052 14272 38108
rect 14272 38052 14328 38108
rect 14328 38052 14332 38108
rect 14268 38048 14332 38052
rect 14348 38108 14412 38112
rect 14348 38052 14352 38108
rect 14352 38052 14408 38108
rect 14408 38052 14412 38108
rect 14348 38048 14412 38052
rect 14428 38108 14492 38112
rect 14428 38052 14432 38108
rect 14432 38052 14488 38108
rect 14488 38052 14492 38108
rect 14428 38048 14492 38052
rect 14508 38108 14572 38112
rect 14508 38052 14512 38108
rect 14512 38052 14568 38108
rect 14568 38052 14572 38108
rect 14508 38048 14572 38052
rect 18707 38108 18771 38112
rect 18707 38052 18711 38108
rect 18711 38052 18767 38108
rect 18767 38052 18771 38108
rect 18707 38048 18771 38052
rect 18787 38108 18851 38112
rect 18787 38052 18791 38108
rect 18791 38052 18847 38108
rect 18847 38052 18851 38108
rect 18787 38048 18851 38052
rect 18867 38108 18931 38112
rect 18867 38052 18871 38108
rect 18871 38052 18927 38108
rect 18927 38052 18931 38108
rect 18867 38048 18931 38052
rect 18947 38108 19011 38112
rect 18947 38052 18951 38108
rect 18951 38052 19007 38108
rect 19007 38052 19011 38108
rect 18947 38048 19011 38052
rect 3171 37564 3235 37568
rect 3171 37508 3175 37564
rect 3175 37508 3231 37564
rect 3231 37508 3235 37564
rect 3171 37504 3235 37508
rect 3251 37564 3315 37568
rect 3251 37508 3255 37564
rect 3255 37508 3311 37564
rect 3311 37508 3315 37564
rect 3251 37504 3315 37508
rect 3331 37564 3395 37568
rect 3331 37508 3335 37564
rect 3335 37508 3391 37564
rect 3391 37508 3395 37564
rect 3331 37504 3395 37508
rect 3411 37564 3475 37568
rect 3411 37508 3415 37564
rect 3415 37508 3471 37564
rect 3471 37508 3475 37564
rect 3411 37504 3475 37508
rect 7610 37564 7674 37568
rect 7610 37508 7614 37564
rect 7614 37508 7670 37564
rect 7670 37508 7674 37564
rect 7610 37504 7674 37508
rect 7690 37564 7754 37568
rect 7690 37508 7694 37564
rect 7694 37508 7750 37564
rect 7750 37508 7754 37564
rect 7690 37504 7754 37508
rect 7770 37564 7834 37568
rect 7770 37508 7774 37564
rect 7774 37508 7830 37564
rect 7830 37508 7834 37564
rect 7770 37504 7834 37508
rect 7850 37564 7914 37568
rect 7850 37508 7854 37564
rect 7854 37508 7910 37564
rect 7910 37508 7914 37564
rect 7850 37504 7914 37508
rect 12049 37564 12113 37568
rect 12049 37508 12053 37564
rect 12053 37508 12109 37564
rect 12109 37508 12113 37564
rect 12049 37504 12113 37508
rect 12129 37564 12193 37568
rect 12129 37508 12133 37564
rect 12133 37508 12189 37564
rect 12189 37508 12193 37564
rect 12129 37504 12193 37508
rect 12209 37564 12273 37568
rect 12209 37508 12213 37564
rect 12213 37508 12269 37564
rect 12269 37508 12273 37564
rect 12209 37504 12273 37508
rect 12289 37564 12353 37568
rect 12289 37508 12293 37564
rect 12293 37508 12349 37564
rect 12349 37508 12353 37564
rect 12289 37504 12353 37508
rect 16488 37564 16552 37568
rect 16488 37508 16492 37564
rect 16492 37508 16548 37564
rect 16548 37508 16552 37564
rect 16488 37504 16552 37508
rect 16568 37564 16632 37568
rect 16568 37508 16572 37564
rect 16572 37508 16628 37564
rect 16628 37508 16632 37564
rect 16568 37504 16632 37508
rect 16648 37564 16712 37568
rect 16648 37508 16652 37564
rect 16652 37508 16708 37564
rect 16708 37508 16712 37564
rect 16648 37504 16712 37508
rect 16728 37564 16792 37568
rect 16728 37508 16732 37564
rect 16732 37508 16788 37564
rect 16788 37508 16792 37564
rect 16728 37504 16792 37508
rect 5390 37020 5454 37024
rect 5390 36964 5394 37020
rect 5394 36964 5450 37020
rect 5450 36964 5454 37020
rect 5390 36960 5454 36964
rect 5470 37020 5534 37024
rect 5470 36964 5474 37020
rect 5474 36964 5530 37020
rect 5530 36964 5534 37020
rect 5470 36960 5534 36964
rect 5550 37020 5614 37024
rect 5550 36964 5554 37020
rect 5554 36964 5610 37020
rect 5610 36964 5614 37020
rect 5550 36960 5614 36964
rect 5630 37020 5694 37024
rect 5630 36964 5634 37020
rect 5634 36964 5690 37020
rect 5690 36964 5694 37020
rect 5630 36960 5694 36964
rect 9829 37020 9893 37024
rect 9829 36964 9833 37020
rect 9833 36964 9889 37020
rect 9889 36964 9893 37020
rect 9829 36960 9893 36964
rect 9909 37020 9973 37024
rect 9909 36964 9913 37020
rect 9913 36964 9969 37020
rect 9969 36964 9973 37020
rect 9909 36960 9973 36964
rect 9989 37020 10053 37024
rect 9989 36964 9993 37020
rect 9993 36964 10049 37020
rect 10049 36964 10053 37020
rect 9989 36960 10053 36964
rect 10069 37020 10133 37024
rect 10069 36964 10073 37020
rect 10073 36964 10129 37020
rect 10129 36964 10133 37020
rect 10069 36960 10133 36964
rect 14268 37020 14332 37024
rect 14268 36964 14272 37020
rect 14272 36964 14328 37020
rect 14328 36964 14332 37020
rect 14268 36960 14332 36964
rect 14348 37020 14412 37024
rect 14348 36964 14352 37020
rect 14352 36964 14408 37020
rect 14408 36964 14412 37020
rect 14348 36960 14412 36964
rect 14428 37020 14492 37024
rect 14428 36964 14432 37020
rect 14432 36964 14488 37020
rect 14488 36964 14492 37020
rect 14428 36960 14492 36964
rect 14508 37020 14572 37024
rect 14508 36964 14512 37020
rect 14512 36964 14568 37020
rect 14568 36964 14572 37020
rect 14508 36960 14572 36964
rect 18707 37020 18771 37024
rect 18707 36964 18711 37020
rect 18711 36964 18767 37020
rect 18767 36964 18771 37020
rect 18707 36960 18771 36964
rect 18787 37020 18851 37024
rect 18787 36964 18791 37020
rect 18791 36964 18847 37020
rect 18847 36964 18851 37020
rect 18787 36960 18851 36964
rect 18867 37020 18931 37024
rect 18867 36964 18871 37020
rect 18871 36964 18927 37020
rect 18927 36964 18931 37020
rect 18867 36960 18931 36964
rect 18947 37020 19011 37024
rect 18947 36964 18951 37020
rect 18951 36964 19007 37020
rect 19007 36964 19011 37020
rect 18947 36960 19011 36964
rect 3171 36476 3235 36480
rect 3171 36420 3175 36476
rect 3175 36420 3231 36476
rect 3231 36420 3235 36476
rect 3171 36416 3235 36420
rect 3251 36476 3315 36480
rect 3251 36420 3255 36476
rect 3255 36420 3311 36476
rect 3311 36420 3315 36476
rect 3251 36416 3315 36420
rect 3331 36476 3395 36480
rect 3331 36420 3335 36476
rect 3335 36420 3391 36476
rect 3391 36420 3395 36476
rect 3331 36416 3395 36420
rect 3411 36476 3475 36480
rect 3411 36420 3415 36476
rect 3415 36420 3471 36476
rect 3471 36420 3475 36476
rect 3411 36416 3475 36420
rect 7610 36476 7674 36480
rect 7610 36420 7614 36476
rect 7614 36420 7670 36476
rect 7670 36420 7674 36476
rect 7610 36416 7674 36420
rect 7690 36476 7754 36480
rect 7690 36420 7694 36476
rect 7694 36420 7750 36476
rect 7750 36420 7754 36476
rect 7690 36416 7754 36420
rect 7770 36476 7834 36480
rect 7770 36420 7774 36476
rect 7774 36420 7830 36476
rect 7830 36420 7834 36476
rect 7770 36416 7834 36420
rect 7850 36476 7914 36480
rect 7850 36420 7854 36476
rect 7854 36420 7910 36476
rect 7910 36420 7914 36476
rect 7850 36416 7914 36420
rect 12049 36476 12113 36480
rect 12049 36420 12053 36476
rect 12053 36420 12109 36476
rect 12109 36420 12113 36476
rect 12049 36416 12113 36420
rect 12129 36476 12193 36480
rect 12129 36420 12133 36476
rect 12133 36420 12189 36476
rect 12189 36420 12193 36476
rect 12129 36416 12193 36420
rect 12209 36476 12273 36480
rect 12209 36420 12213 36476
rect 12213 36420 12269 36476
rect 12269 36420 12273 36476
rect 12209 36416 12273 36420
rect 12289 36476 12353 36480
rect 12289 36420 12293 36476
rect 12293 36420 12349 36476
rect 12349 36420 12353 36476
rect 12289 36416 12353 36420
rect 16488 36476 16552 36480
rect 16488 36420 16492 36476
rect 16492 36420 16548 36476
rect 16548 36420 16552 36476
rect 16488 36416 16552 36420
rect 16568 36476 16632 36480
rect 16568 36420 16572 36476
rect 16572 36420 16628 36476
rect 16628 36420 16632 36476
rect 16568 36416 16632 36420
rect 16648 36476 16712 36480
rect 16648 36420 16652 36476
rect 16652 36420 16708 36476
rect 16708 36420 16712 36476
rect 16648 36416 16712 36420
rect 16728 36476 16792 36480
rect 16728 36420 16732 36476
rect 16732 36420 16788 36476
rect 16788 36420 16792 36476
rect 16728 36416 16792 36420
rect 5390 35932 5454 35936
rect 5390 35876 5394 35932
rect 5394 35876 5450 35932
rect 5450 35876 5454 35932
rect 5390 35872 5454 35876
rect 5470 35932 5534 35936
rect 5470 35876 5474 35932
rect 5474 35876 5530 35932
rect 5530 35876 5534 35932
rect 5470 35872 5534 35876
rect 5550 35932 5614 35936
rect 5550 35876 5554 35932
rect 5554 35876 5610 35932
rect 5610 35876 5614 35932
rect 5550 35872 5614 35876
rect 5630 35932 5694 35936
rect 5630 35876 5634 35932
rect 5634 35876 5690 35932
rect 5690 35876 5694 35932
rect 5630 35872 5694 35876
rect 9829 35932 9893 35936
rect 9829 35876 9833 35932
rect 9833 35876 9889 35932
rect 9889 35876 9893 35932
rect 9829 35872 9893 35876
rect 9909 35932 9973 35936
rect 9909 35876 9913 35932
rect 9913 35876 9969 35932
rect 9969 35876 9973 35932
rect 9909 35872 9973 35876
rect 9989 35932 10053 35936
rect 9989 35876 9993 35932
rect 9993 35876 10049 35932
rect 10049 35876 10053 35932
rect 9989 35872 10053 35876
rect 10069 35932 10133 35936
rect 10069 35876 10073 35932
rect 10073 35876 10129 35932
rect 10129 35876 10133 35932
rect 10069 35872 10133 35876
rect 14268 35932 14332 35936
rect 14268 35876 14272 35932
rect 14272 35876 14328 35932
rect 14328 35876 14332 35932
rect 14268 35872 14332 35876
rect 14348 35932 14412 35936
rect 14348 35876 14352 35932
rect 14352 35876 14408 35932
rect 14408 35876 14412 35932
rect 14348 35872 14412 35876
rect 14428 35932 14492 35936
rect 14428 35876 14432 35932
rect 14432 35876 14488 35932
rect 14488 35876 14492 35932
rect 14428 35872 14492 35876
rect 14508 35932 14572 35936
rect 14508 35876 14512 35932
rect 14512 35876 14568 35932
rect 14568 35876 14572 35932
rect 14508 35872 14572 35876
rect 18707 35932 18771 35936
rect 18707 35876 18711 35932
rect 18711 35876 18767 35932
rect 18767 35876 18771 35932
rect 18707 35872 18771 35876
rect 18787 35932 18851 35936
rect 18787 35876 18791 35932
rect 18791 35876 18847 35932
rect 18847 35876 18851 35932
rect 18787 35872 18851 35876
rect 18867 35932 18931 35936
rect 18867 35876 18871 35932
rect 18871 35876 18927 35932
rect 18927 35876 18931 35932
rect 18867 35872 18931 35876
rect 18947 35932 19011 35936
rect 18947 35876 18951 35932
rect 18951 35876 19007 35932
rect 19007 35876 19011 35932
rect 18947 35872 19011 35876
rect 3171 35388 3235 35392
rect 3171 35332 3175 35388
rect 3175 35332 3231 35388
rect 3231 35332 3235 35388
rect 3171 35328 3235 35332
rect 3251 35388 3315 35392
rect 3251 35332 3255 35388
rect 3255 35332 3311 35388
rect 3311 35332 3315 35388
rect 3251 35328 3315 35332
rect 3331 35388 3395 35392
rect 3331 35332 3335 35388
rect 3335 35332 3391 35388
rect 3391 35332 3395 35388
rect 3331 35328 3395 35332
rect 3411 35388 3475 35392
rect 3411 35332 3415 35388
rect 3415 35332 3471 35388
rect 3471 35332 3475 35388
rect 3411 35328 3475 35332
rect 7610 35388 7674 35392
rect 7610 35332 7614 35388
rect 7614 35332 7670 35388
rect 7670 35332 7674 35388
rect 7610 35328 7674 35332
rect 7690 35388 7754 35392
rect 7690 35332 7694 35388
rect 7694 35332 7750 35388
rect 7750 35332 7754 35388
rect 7690 35328 7754 35332
rect 7770 35388 7834 35392
rect 7770 35332 7774 35388
rect 7774 35332 7830 35388
rect 7830 35332 7834 35388
rect 7770 35328 7834 35332
rect 7850 35388 7914 35392
rect 7850 35332 7854 35388
rect 7854 35332 7910 35388
rect 7910 35332 7914 35388
rect 7850 35328 7914 35332
rect 12049 35388 12113 35392
rect 12049 35332 12053 35388
rect 12053 35332 12109 35388
rect 12109 35332 12113 35388
rect 12049 35328 12113 35332
rect 12129 35388 12193 35392
rect 12129 35332 12133 35388
rect 12133 35332 12189 35388
rect 12189 35332 12193 35388
rect 12129 35328 12193 35332
rect 12209 35388 12273 35392
rect 12209 35332 12213 35388
rect 12213 35332 12269 35388
rect 12269 35332 12273 35388
rect 12209 35328 12273 35332
rect 12289 35388 12353 35392
rect 12289 35332 12293 35388
rect 12293 35332 12349 35388
rect 12349 35332 12353 35388
rect 12289 35328 12353 35332
rect 16488 35388 16552 35392
rect 16488 35332 16492 35388
rect 16492 35332 16548 35388
rect 16548 35332 16552 35388
rect 16488 35328 16552 35332
rect 16568 35388 16632 35392
rect 16568 35332 16572 35388
rect 16572 35332 16628 35388
rect 16628 35332 16632 35388
rect 16568 35328 16632 35332
rect 16648 35388 16712 35392
rect 16648 35332 16652 35388
rect 16652 35332 16708 35388
rect 16708 35332 16712 35388
rect 16648 35328 16712 35332
rect 16728 35388 16792 35392
rect 16728 35332 16732 35388
rect 16732 35332 16788 35388
rect 16788 35332 16792 35388
rect 16728 35328 16792 35332
rect 5390 34844 5454 34848
rect 5390 34788 5394 34844
rect 5394 34788 5450 34844
rect 5450 34788 5454 34844
rect 5390 34784 5454 34788
rect 5470 34844 5534 34848
rect 5470 34788 5474 34844
rect 5474 34788 5530 34844
rect 5530 34788 5534 34844
rect 5470 34784 5534 34788
rect 5550 34844 5614 34848
rect 5550 34788 5554 34844
rect 5554 34788 5610 34844
rect 5610 34788 5614 34844
rect 5550 34784 5614 34788
rect 5630 34844 5694 34848
rect 5630 34788 5634 34844
rect 5634 34788 5690 34844
rect 5690 34788 5694 34844
rect 5630 34784 5694 34788
rect 9829 34844 9893 34848
rect 9829 34788 9833 34844
rect 9833 34788 9889 34844
rect 9889 34788 9893 34844
rect 9829 34784 9893 34788
rect 9909 34844 9973 34848
rect 9909 34788 9913 34844
rect 9913 34788 9969 34844
rect 9969 34788 9973 34844
rect 9909 34784 9973 34788
rect 9989 34844 10053 34848
rect 9989 34788 9993 34844
rect 9993 34788 10049 34844
rect 10049 34788 10053 34844
rect 9989 34784 10053 34788
rect 10069 34844 10133 34848
rect 10069 34788 10073 34844
rect 10073 34788 10129 34844
rect 10129 34788 10133 34844
rect 10069 34784 10133 34788
rect 14268 34844 14332 34848
rect 14268 34788 14272 34844
rect 14272 34788 14328 34844
rect 14328 34788 14332 34844
rect 14268 34784 14332 34788
rect 14348 34844 14412 34848
rect 14348 34788 14352 34844
rect 14352 34788 14408 34844
rect 14408 34788 14412 34844
rect 14348 34784 14412 34788
rect 14428 34844 14492 34848
rect 14428 34788 14432 34844
rect 14432 34788 14488 34844
rect 14488 34788 14492 34844
rect 14428 34784 14492 34788
rect 14508 34844 14572 34848
rect 14508 34788 14512 34844
rect 14512 34788 14568 34844
rect 14568 34788 14572 34844
rect 14508 34784 14572 34788
rect 18707 34844 18771 34848
rect 18707 34788 18711 34844
rect 18711 34788 18767 34844
rect 18767 34788 18771 34844
rect 18707 34784 18771 34788
rect 18787 34844 18851 34848
rect 18787 34788 18791 34844
rect 18791 34788 18847 34844
rect 18847 34788 18851 34844
rect 18787 34784 18851 34788
rect 18867 34844 18931 34848
rect 18867 34788 18871 34844
rect 18871 34788 18927 34844
rect 18927 34788 18931 34844
rect 18867 34784 18931 34788
rect 18947 34844 19011 34848
rect 18947 34788 18951 34844
rect 18951 34788 19007 34844
rect 19007 34788 19011 34844
rect 18947 34784 19011 34788
rect 3171 34300 3235 34304
rect 3171 34244 3175 34300
rect 3175 34244 3231 34300
rect 3231 34244 3235 34300
rect 3171 34240 3235 34244
rect 3251 34300 3315 34304
rect 3251 34244 3255 34300
rect 3255 34244 3311 34300
rect 3311 34244 3315 34300
rect 3251 34240 3315 34244
rect 3331 34300 3395 34304
rect 3331 34244 3335 34300
rect 3335 34244 3391 34300
rect 3391 34244 3395 34300
rect 3331 34240 3395 34244
rect 3411 34300 3475 34304
rect 3411 34244 3415 34300
rect 3415 34244 3471 34300
rect 3471 34244 3475 34300
rect 3411 34240 3475 34244
rect 7610 34300 7674 34304
rect 7610 34244 7614 34300
rect 7614 34244 7670 34300
rect 7670 34244 7674 34300
rect 7610 34240 7674 34244
rect 7690 34300 7754 34304
rect 7690 34244 7694 34300
rect 7694 34244 7750 34300
rect 7750 34244 7754 34300
rect 7690 34240 7754 34244
rect 7770 34300 7834 34304
rect 7770 34244 7774 34300
rect 7774 34244 7830 34300
rect 7830 34244 7834 34300
rect 7770 34240 7834 34244
rect 7850 34300 7914 34304
rect 7850 34244 7854 34300
rect 7854 34244 7910 34300
rect 7910 34244 7914 34300
rect 7850 34240 7914 34244
rect 12049 34300 12113 34304
rect 12049 34244 12053 34300
rect 12053 34244 12109 34300
rect 12109 34244 12113 34300
rect 12049 34240 12113 34244
rect 12129 34300 12193 34304
rect 12129 34244 12133 34300
rect 12133 34244 12189 34300
rect 12189 34244 12193 34300
rect 12129 34240 12193 34244
rect 12209 34300 12273 34304
rect 12209 34244 12213 34300
rect 12213 34244 12269 34300
rect 12269 34244 12273 34300
rect 12209 34240 12273 34244
rect 12289 34300 12353 34304
rect 12289 34244 12293 34300
rect 12293 34244 12349 34300
rect 12349 34244 12353 34300
rect 12289 34240 12353 34244
rect 16488 34300 16552 34304
rect 16488 34244 16492 34300
rect 16492 34244 16548 34300
rect 16548 34244 16552 34300
rect 16488 34240 16552 34244
rect 16568 34300 16632 34304
rect 16568 34244 16572 34300
rect 16572 34244 16628 34300
rect 16628 34244 16632 34300
rect 16568 34240 16632 34244
rect 16648 34300 16712 34304
rect 16648 34244 16652 34300
rect 16652 34244 16708 34300
rect 16708 34244 16712 34300
rect 16648 34240 16712 34244
rect 16728 34300 16792 34304
rect 16728 34244 16732 34300
rect 16732 34244 16788 34300
rect 16788 34244 16792 34300
rect 16728 34240 16792 34244
rect 5390 33756 5454 33760
rect 5390 33700 5394 33756
rect 5394 33700 5450 33756
rect 5450 33700 5454 33756
rect 5390 33696 5454 33700
rect 5470 33756 5534 33760
rect 5470 33700 5474 33756
rect 5474 33700 5530 33756
rect 5530 33700 5534 33756
rect 5470 33696 5534 33700
rect 5550 33756 5614 33760
rect 5550 33700 5554 33756
rect 5554 33700 5610 33756
rect 5610 33700 5614 33756
rect 5550 33696 5614 33700
rect 5630 33756 5694 33760
rect 5630 33700 5634 33756
rect 5634 33700 5690 33756
rect 5690 33700 5694 33756
rect 5630 33696 5694 33700
rect 9829 33756 9893 33760
rect 9829 33700 9833 33756
rect 9833 33700 9889 33756
rect 9889 33700 9893 33756
rect 9829 33696 9893 33700
rect 9909 33756 9973 33760
rect 9909 33700 9913 33756
rect 9913 33700 9969 33756
rect 9969 33700 9973 33756
rect 9909 33696 9973 33700
rect 9989 33756 10053 33760
rect 9989 33700 9993 33756
rect 9993 33700 10049 33756
rect 10049 33700 10053 33756
rect 9989 33696 10053 33700
rect 10069 33756 10133 33760
rect 10069 33700 10073 33756
rect 10073 33700 10129 33756
rect 10129 33700 10133 33756
rect 10069 33696 10133 33700
rect 14268 33756 14332 33760
rect 14268 33700 14272 33756
rect 14272 33700 14328 33756
rect 14328 33700 14332 33756
rect 14268 33696 14332 33700
rect 14348 33756 14412 33760
rect 14348 33700 14352 33756
rect 14352 33700 14408 33756
rect 14408 33700 14412 33756
rect 14348 33696 14412 33700
rect 14428 33756 14492 33760
rect 14428 33700 14432 33756
rect 14432 33700 14488 33756
rect 14488 33700 14492 33756
rect 14428 33696 14492 33700
rect 14508 33756 14572 33760
rect 14508 33700 14512 33756
rect 14512 33700 14568 33756
rect 14568 33700 14572 33756
rect 14508 33696 14572 33700
rect 18707 33756 18771 33760
rect 18707 33700 18711 33756
rect 18711 33700 18767 33756
rect 18767 33700 18771 33756
rect 18707 33696 18771 33700
rect 18787 33756 18851 33760
rect 18787 33700 18791 33756
rect 18791 33700 18847 33756
rect 18847 33700 18851 33756
rect 18787 33696 18851 33700
rect 18867 33756 18931 33760
rect 18867 33700 18871 33756
rect 18871 33700 18927 33756
rect 18927 33700 18931 33756
rect 18867 33696 18931 33700
rect 18947 33756 19011 33760
rect 18947 33700 18951 33756
rect 18951 33700 19007 33756
rect 19007 33700 19011 33756
rect 18947 33696 19011 33700
rect 3171 33212 3235 33216
rect 3171 33156 3175 33212
rect 3175 33156 3231 33212
rect 3231 33156 3235 33212
rect 3171 33152 3235 33156
rect 3251 33212 3315 33216
rect 3251 33156 3255 33212
rect 3255 33156 3311 33212
rect 3311 33156 3315 33212
rect 3251 33152 3315 33156
rect 3331 33212 3395 33216
rect 3331 33156 3335 33212
rect 3335 33156 3391 33212
rect 3391 33156 3395 33212
rect 3331 33152 3395 33156
rect 3411 33212 3475 33216
rect 3411 33156 3415 33212
rect 3415 33156 3471 33212
rect 3471 33156 3475 33212
rect 3411 33152 3475 33156
rect 7610 33212 7674 33216
rect 7610 33156 7614 33212
rect 7614 33156 7670 33212
rect 7670 33156 7674 33212
rect 7610 33152 7674 33156
rect 7690 33212 7754 33216
rect 7690 33156 7694 33212
rect 7694 33156 7750 33212
rect 7750 33156 7754 33212
rect 7690 33152 7754 33156
rect 7770 33212 7834 33216
rect 7770 33156 7774 33212
rect 7774 33156 7830 33212
rect 7830 33156 7834 33212
rect 7770 33152 7834 33156
rect 7850 33212 7914 33216
rect 7850 33156 7854 33212
rect 7854 33156 7910 33212
rect 7910 33156 7914 33212
rect 7850 33152 7914 33156
rect 12049 33212 12113 33216
rect 12049 33156 12053 33212
rect 12053 33156 12109 33212
rect 12109 33156 12113 33212
rect 12049 33152 12113 33156
rect 12129 33212 12193 33216
rect 12129 33156 12133 33212
rect 12133 33156 12189 33212
rect 12189 33156 12193 33212
rect 12129 33152 12193 33156
rect 12209 33212 12273 33216
rect 12209 33156 12213 33212
rect 12213 33156 12269 33212
rect 12269 33156 12273 33212
rect 12209 33152 12273 33156
rect 12289 33212 12353 33216
rect 12289 33156 12293 33212
rect 12293 33156 12349 33212
rect 12349 33156 12353 33212
rect 12289 33152 12353 33156
rect 16488 33212 16552 33216
rect 16488 33156 16492 33212
rect 16492 33156 16548 33212
rect 16548 33156 16552 33212
rect 16488 33152 16552 33156
rect 16568 33212 16632 33216
rect 16568 33156 16572 33212
rect 16572 33156 16628 33212
rect 16628 33156 16632 33212
rect 16568 33152 16632 33156
rect 16648 33212 16712 33216
rect 16648 33156 16652 33212
rect 16652 33156 16708 33212
rect 16708 33156 16712 33212
rect 16648 33152 16712 33156
rect 16728 33212 16792 33216
rect 16728 33156 16732 33212
rect 16732 33156 16788 33212
rect 16788 33156 16792 33212
rect 16728 33152 16792 33156
rect 5390 32668 5454 32672
rect 5390 32612 5394 32668
rect 5394 32612 5450 32668
rect 5450 32612 5454 32668
rect 5390 32608 5454 32612
rect 5470 32668 5534 32672
rect 5470 32612 5474 32668
rect 5474 32612 5530 32668
rect 5530 32612 5534 32668
rect 5470 32608 5534 32612
rect 5550 32668 5614 32672
rect 5550 32612 5554 32668
rect 5554 32612 5610 32668
rect 5610 32612 5614 32668
rect 5550 32608 5614 32612
rect 5630 32668 5694 32672
rect 5630 32612 5634 32668
rect 5634 32612 5690 32668
rect 5690 32612 5694 32668
rect 5630 32608 5694 32612
rect 9829 32668 9893 32672
rect 9829 32612 9833 32668
rect 9833 32612 9889 32668
rect 9889 32612 9893 32668
rect 9829 32608 9893 32612
rect 9909 32668 9973 32672
rect 9909 32612 9913 32668
rect 9913 32612 9969 32668
rect 9969 32612 9973 32668
rect 9909 32608 9973 32612
rect 9989 32668 10053 32672
rect 9989 32612 9993 32668
rect 9993 32612 10049 32668
rect 10049 32612 10053 32668
rect 9989 32608 10053 32612
rect 10069 32668 10133 32672
rect 10069 32612 10073 32668
rect 10073 32612 10129 32668
rect 10129 32612 10133 32668
rect 10069 32608 10133 32612
rect 14268 32668 14332 32672
rect 14268 32612 14272 32668
rect 14272 32612 14328 32668
rect 14328 32612 14332 32668
rect 14268 32608 14332 32612
rect 14348 32668 14412 32672
rect 14348 32612 14352 32668
rect 14352 32612 14408 32668
rect 14408 32612 14412 32668
rect 14348 32608 14412 32612
rect 14428 32668 14492 32672
rect 14428 32612 14432 32668
rect 14432 32612 14488 32668
rect 14488 32612 14492 32668
rect 14428 32608 14492 32612
rect 14508 32668 14572 32672
rect 14508 32612 14512 32668
rect 14512 32612 14568 32668
rect 14568 32612 14572 32668
rect 14508 32608 14572 32612
rect 18707 32668 18771 32672
rect 18707 32612 18711 32668
rect 18711 32612 18767 32668
rect 18767 32612 18771 32668
rect 18707 32608 18771 32612
rect 18787 32668 18851 32672
rect 18787 32612 18791 32668
rect 18791 32612 18847 32668
rect 18847 32612 18851 32668
rect 18787 32608 18851 32612
rect 18867 32668 18931 32672
rect 18867 32612 18871 32668
rect 18871 32612 18927 32668
rect 18927 32612 18931 32668
rect 18867 32608 18931 32612
rect 18947 32668 19011 32672
rect 18947 32612 18951 32668
rect 18951 32612 19007 32668
rect 19007 32612 19011 32668
rect 18947 32608 19011 32612
rect 3171 32124 3235 32128
rect 3171 32068 3175 32124
rect 3175 32068 3231 32124
rect 3231 32068 3235 32124
rect 3171 32064 3235 32068
rect 3251 32124 3315 32128
rect 3251 32068 3255 32124
rect 3255 32068 3311 32124
rect 3311 32068 3315 32124
rect 3251 32064 3315 32068
rect 3331 32124 3395 32128
rect 3331 32068 3335 32124
rect 3335 32068 3391 32124
rect 3391 32068 3395 32124
rect 3331 32064 3395 32068
rect 3411 32124 3475 32128
rect 3411 32068 3415 32124
rect 3415 32068 3471 32124
rect 3471 32068 3475 32124
rect 3411 32064 3475 32068
rect 7610 32124 7674 32128
rect 7610 32068 7614 32124
rect 7614 32068 7670 32124
rect 7670 32068 7674 32124
rect 7610 32064 7674 32068
rect 7690 32124 7754 32128
rect 7690 32068 7694 32124
rect 7694 32068 7750 32124
rect 7750 32068 7754 32124
rect 7690 32064 7754 32068
rect 7770 32124 7834 32128
rect 7770 32068 7774 32124
rect 7774 32068 7830 32124
rect 7830 32068 7834 32124
rect 7770 32064 7834 32068
rect 7850 32124 7914 32128
rect 7850 32068 7854 32124
rect 7854 32068 7910 32124
rect 7910 32068 7914 32124
rect 7850 32064 7914 32068
rect 12049 32124 12113 32128
rect 12049 32068 12053 32124
rect 12053 32068 12109 32124
rect 12109 32068 12113 32124
rect 12049 32064 12113 32068
rect 12129 32124 12193 32128
rect 12129 32068 12133 32124
rect 12133 32068 12189 32124
rect 12189 32068 12193 32124
rect 12129 32064 12193 32068
rect 12209 32124 12273 32128
rect 12209 32068 12213 32124
rect 12213 32068 12269 32124
rect 12269 32068 12273 32124
rect 12209 32064 12273 32068
rect 12289 32124 12353 32128
rect 12289 32068 12293 32124
rect 12293 32068 12349 32124
rect 12349 32068 12353 32124
rect 12289 32064 12353 32068
rect 16488 32124 16552 32128
rect 16488 32068 16492 32124
rect 16492 32068 16548 32124
rect 16548 32068 16552 32124
rect 16488 32064 16552 32068
rect 16568 32124 16632 32128
rect 16568 32068 16572 32124
rect 16572 32068 16628 32124
rect 16628 32068 16632 32124
rect 16568 32064 16632 32068
rect 16648 32124 16712 32128
rect 16648 32068 16652 32124
rect 16652 32068 16708 32124
rect 16708 32068 16712 32124
rect 16648 32064 16712 32068
rect 16728 32124 16792 32128
rect 16728 32068 16732 32124
rect 16732 32068 16788 32124
rect 16788 32068 16792 32124
rect 16728 32064 16792 32068
rect 5390 31580 5454 31584
rect 5390 31524 5394 31580
rect 5394 31524 5450 31580
rect 5450 31524 5454 31580
rect 5390 31520 5454 31524
rect 5470 31580 5534 31584
rect 5470 31524 5474 31580
rect 5474 31524 5530 31580
rect 5530 31524 5534 31580
rect 5470 31520 5534 31524
rect 5550 31580 5614 31584
rect 5550 31524 5554 31580
rect 5554 31524 5610 31580
rect 5610 31524 5614 31580
rect 5550 31520 5614 31524
rect 5630 31580 5694 31584
rect 5630 31524 5634 31580
rect 5634 31524 5690 31580
rect 5690 31524 5694 31580
rect 5630 31520 5694 31524
rect 9829 31580 9893 31584
rect 9829 31524 9833 31580
rect 9833 31524 9889 31580
rect 9889 31524 9893 31580
rect 9829 31520 9893 31524
rect 9909 31580 9973 31584
rect 9909 31524 9913 31580
rect 9913 31524 9969 31580
rect 9969 31524 9973 31580
rect 9909 31520 9973 31524
rect 9989 31580 10053 31584
rect 9989 31524 9993 31580
rect 9993 31524 10049 31580
rect 10049 31524 10053 31580
rect 9989 31520 10053 31524
rect 10069 31580 10133 31584
rect 10069 31524 10073 31580
rect 10073 31524 10129 31580
rect 10129 31524 10133 31580
rect 10069 31520 10133 31524
rect 14268 31580 14332 31584
rect 14268 31524 14272 31580
rect 14272 31524 14328 31580
rect 14328 31524 14332 31580
rect 14268 31520 14332 31524
rect 14348 31580 14412 31584
rect 14348 31524 14352 31580
rect 14352 31524 14408 31580
rect 14408 31524 14412 31580
rect 14348 31520 14412 31524
rect 14428 31580 14492 31584
rect 14428 31524 14432 31580
rect 14432 31524 14488 31580
rect 14488 31524 14492 31580
rect 14428 31520 14492 31524
rect 14508 31580 14572 31584
rect 14508 31524 14512 31580
rect 14512 31524 14568 31580
rect 14568 31524 14572 31580
rect 14508 31520 14572 31524
rect 18707 31580 18771 31584
rect 18707 31524 18711 31580
rect 18711 31524 18767 31580
rect 18767 31524 18771 31580
rect 18707 31520 18771 31524
rect 18787 31580 18851 31584
rect 18787 31524 18791 31580
rect 18791 31524 18847 31580
rect 18847 31524 18851 31580
rect 18787 31520 18851 31524
rect 18867 31580 18931 31584
rect 18867 31524 18871 31580
rect 18871 31524 18927 31580
rect 18927 31524 18931 31580
rect 18867 31520 18931 31524
rect 18947 31580 19011 31584
rect 18947 31524 18951 31580
rect 18951 31524 19007 31580
rect 19007 31524 19011 31580
rect 18947 31520 19011 31524
rect 3171 31036 3235 31040
rect 3171 30980 3175 31036
rect 3175 30980 3231 31036
rect 3231 30980 3235 31036
rect 3171 30976 3235 30980
rect 3251 31036 3315 31040
rect 3251 30980 3255 31036
rect 3255 30980 3311 31036
rect 3311 30980 3315 31036
rect 3251 30976 3315 30980
rect 3331 31036 3395 31040
rect 3331 30980 3335 31036
rect 3335 30980 3391 31036
rect 3391 30980 3395 31036
rect 3331 30976 3395 30980
rect 3411 31036 3475 31040
rect 3411 30980 3415 31036
rect 3415 30980 3471 31036
rect 3471 30980 3475 31036
rect 3411 30976 3475 30980
rect 7610 31036 7674 31040
rect 7610 30980 7614 31036
rect 7614 30980 7670 31036
rect 7670 30980 7674 31036
rect 7610 30976 7674 30980
rect 7690 31036 7754 31040
rect 7690 30980 7694 31036
rect 7694 30980 7750 31036
rect 7750 30980 7754 31036
rect 7690 30976 7754 30980
rect 7770 31036 7834 31040
rect 7770 30980 7774 31036
rect 7774 30980 7830 31036
rect 7830 30980 7834 31036
rect 7770 30976 7834 30980
rect 7850 31036 7914 31040
rect 7850 30980 7854 31036
rect 7854 30980 7910 31036
rect 7910 30980 7914 31036
rect 7850 30976 7914 30980
rect 12049 31036 12113 31040
rect 12049 30980 12053 31036
rect 12053 30980 12109 31036
rect 12109 30980 12113 31036
rect 12049 30976 12113 30980
rect 12129 31036 12193 31040
rect 12129 30980 12133 31036
rect 12133 30980 12189 31036
rect 12189 30980 12193 31036
rect 12129 30976 12193 30980
rect 12209 31036 12273 31040
rect 12209 30980 12213 31036
rect 12213 30980 12269 31036
rect 12269 30980 12273 31036
rect 12209 30976 12273 30980
rect 12289 31036 12353 31040
rect 12289 30980 12293 31036
rect 12293 30980 12349 31036
rect 12349 30980 12353 31036
rect 12289 30976 12353 30980
rect 16488 31036 16552 31040
rect 16488 30980 16492 31036
rect 16492 30980 16548 31036
rect 16548 30980 16552 31036
rect 16488 30976 16552 30980
rect 16568 31036 16632 31040
rect 16568 30980 16572 31036
rect 16572 30980 16628 31036
rect 16628 30980 16632 31036
rect 16568 30976 16632 30980
rect 16648 31036 16712 31040
rect 16648 30980 16652 31036
rect 16652 30980 16708 31036
rect 16708 30980 16712 31036
rect 16648 30976 16712 30980
rect 16728 31036 16792 31040
rect 16728 30980 16732 31036
rect 16732 30980 16788 31036
rect 16788 30980 16792 31036
rect 16728 30976 16792 30980
rect 5390 30492 5454 30496
rect 5390 30436 5394 30492
rect 5394 30436 5450 30492
rect 5450 30436 5454 30492
rect 5390 30432 5454 30436
rect 5470 30492 5534 30496
rect 5470 30436 5474 30492
rect 5474 30436 5530 30492
rect 5530 30436 5534 30492
rect 5470 30432 5534 30436
rect 5550 30492 5614 30496
rect 5550 30436 5554 30492
rect 5554 30436 5610 30492
rect 5610 30436 5614 30492
rect 5550 30432 5614 30436
rect 5630 30492 5694 30496
rect 5630 30436 5634 30492
rect 5634 30436 5690 30492
rect 5690 30436 5694 30492
rect 5630 30432 5694 30436
rect 9829 30492 9893 30496
rect 9829 30436 9833 30492
rect 9833 30436 9889 30492
rect 9889 30436 9893 30492
rect 9829 30432 9893 30436
rect 9909 30492 9973 30496
rect 9909 30436 9913 30492
rect 9913 30436 9969 30492
rect 9969 30436 9973 30492
rect 9909 30432 9973 30436
rect 9989 30492 10053 30496
rect 9989 30436 9993 30492
rect 9993 30436 10049 30492
rect 10049 30436 10053 30492
rect 9989 30432 10053 30436
rect 10069 30492 10133 30496
rect 10069 30436 10073 30492
rect 10073 30436 10129 30492
rect 10129 30436 10133 30492
rect 10069 30432 10133 30436
rect 14268 30492 14332 30496
rect 14268 30436 14272 30492
rect 14272 30436 14328 30492
rect 14328 30436 14332 30492
rect 14268 30432 14332 30436
rect 14348 30492 14412 30496
rect 14348 30436 14352 30492
rect 14352 30436 14408 30492
rect 14408 30436 14412 30492
rect 14348 30432 14412 30436
rect 14428 30492 14492 30496
rect 14428 30436 14432 30492
rect 14432 30436 14488 30492
rect 14488 30436 14492 30492
rect 14428 30432 14492 30436
rect 14508 30492 14572 30496
rect 14508 30436 14512 30492
rect 14512 30436 14568 30492
rect 14568 30436 14572 30492
rect 14508 30432 14572 30436
rect 18707 30492 18771 30496
rect 18707 30436 18711 30492
rect 18711 30436 18767 30492
rect 18767 30436 18771 30492
rect 18707 30432 18771 30436
rect 18787 30492 18851 30496
rect 18787 30436 18791 30492
rect 18791 30436 18847 30492
rect 18847 30436 18851 30492
rect 18787 30432 18851 30436
rect 18867 30492 18931 30496
rect 18867 30436 18871 30492
rect 18871 30436 18927 30492
rect 18927 30436 18931 30492
rect 18867 30432 18931 30436
rect 18947 30492 19011 30496
rect 18947 30436 18951 30492
rect 18951 30436 19007 30492
rect 19007 30436 19011 30492
rect 18947 30432 19011 30436
rect 3171 29948 3235 29952
rect 3171 29892 3175 29948
rect 3175 29892 3231 29948
rect 3231 29892 3235 29948
rect 3171 29888 3235 29892
rect 3251 29948 3315 29952
rect 3251 29892 3255 29948
rect 3255 29892 3311 29948
rect 3311 29892 3315 29948
rect 3251 29888 3315 29892
rect 3331 29948 3395 29952
rect 3331 29892 3335 29948
rect 3335 29892 3391 29948
rect 3391 29892 3395 29948
rect 3331 29888 3395 29892
rect 3411 29948 3475 29952
rect 3411 29892 3415 29948
rect 3415 29892 3471 29948
rect 3471 29892 3475 29948
rect 3411 29888 3475 29892
rect 7610 29948 7674 29952
rect 7610 29892 7614 29948
rect 7614 29892 7670 29948
rect 7670 29892 7674 29948
rect 7610 29888 7674 29892
rect 7690 29948 7754 29952
rect 7690 29892 7694 29948
rect 7694 29892 7750 29948
rect 7750 29892 7754 29948
rect 7690 29888 7754 29892
rect 7770 29948 7834 29952
rect 7770 29892 7774 29948
rect 7774 29892 7830 29948
rect 7830 29892 7834 29948
rect 7770 29888 7834 29892
rect 7850 29948 7914 29952
rect 7850 29892 7854 29948
rect 7854 29892 7910 29948
rect 7910 29892 7914 29948
rect 7850 29888 7914 29892
rect 12049 29948 12113 29952
rect 12049 29892 12053 29948
rect 12053 29892 12109 29948
rect 12109 29892 12113 29948
rect 12049 29888 12113 29892
rect 12129 29948 12193 29952
rect 12129 29892 12133 29948
rect 12133 29892 12189 29948
rect 12189 29892 12193 29948
rect 12129 29888 12193 29892
rect 12209 29948 12273 29952
rect 12209 29892 12213 29948
rect 12213 29892 12269 29948
rect 12269 29892 12273 29948
rect 12209 29888 12273 29892
rect 12289 29948 12353 29952
rect 12289 29892 12293 29948
rect 12293 29892 12349 29948
rect 12349 29892 12353 29948
rect 12289 29888 12353 29892
rect 16488 29948 16552 29952
rect 16488 29892 16492 29948
rect 16492 29892 16548 29948
rect 16548 29892 16552 29948
rect 16488 29888 16552 29892
rect 16568 29948 16632 29952
rect 16568 29892 16572 29948
rect 16572 29892 16628 29948
rect 16628 29892 16632 29948
rect 16568 29888 16632 29892
rect 16648 29948 16712 29952
rect 16648 29892 16652 29948
rect 16652 29892 16708 29948
rect 16708 29892 16712 29948
rect 16648 29888 16712 29892
rect 16728 29948 16792 29952
rect 16728 29892 16732 29948
rect 16732 29892 16788 29948
rect 16788 29892 16792 29948
rect 16728 29888 16792 29892
rect 5390 29404 5454 29408
rect 5390 29348 5394 29404
rect 5394 29348 5450 29404
rect 5450 29348 5454 29404
rect 5390 29344 5454 29348
rect 5470 29404 5534 29408
rect 5470 29348 5474 29404
rect 5474 29348 5530 29404
rect 5530 29348 5534 29404
rect 5470 29344 5534 29348
rect 5550 29404 5614 29408
rect 5550 29348 5554 29404
rect 5554 29348 5610 29404
rect 5610 29348 5614 29404
rect 5550 29344 5614 29348
rect 5630 29404 5694 29408
rect 5630 29348 5634 29404
rect 5634 29348 5690 29404
rect 5690 29348 5694 29404
rect 5630 29344 5694 29348
rect 9829 29404 9893 29408
rect 9829 29348 9833 29404
rect 9833 29348 9889 29404
rect 9889 29348 9893 29404
rect 9829 29344 9893 29348
rect 9909 29404 9973 29408
rect 9909 29348 9913 29404
rect 9913 29348 9969 29404
rect 9969 29348 9973 29404
rect 9909 29344 9973 29348
rect 9989 29404 10053 29408
rect 9989 29348 9993 29404
rect 9993 29348 10049 29404
rect 10049 29348 10053 29404
rect 9989 29344 10053 29348
rect 10069 29404 10133 29408
rect 10069 29348 10073 29404
rect 10073 29348 10129 29404
rect 10129 29348 10133 29404
rect 10069 29344 10133 29348
rect 14268 29404 14332 29408
rect 14268 29348 14272 29404
rect 14272 29348 14328 29404
rect 14328 29348 14332 29404
rect 14268 29344 14332 29348
rect 14348 29404 14412 29408
rect 14348 29348 14352 29404
rect 14352 29348 14408 29404
rect 14408 29348 14412 29404
rect 14348 29344 14412 29348
rect 14428 29404 14492 29408
rect 14428 29348 14432 29404
rect 14432 29348 14488 29404
rect 14488 29348 14492 29404
rect 14428 29344 14492 29348
rect 14508 29404 14572 29408
rect 14508 29348 14512 29404
rect 14512 29348 14568 29404
rect 14568 29348 14572 29404
rect 14508 29344 14572 29348
rect 18707 29404 18771 29408
rect 18707 29348 18711 29404
rect 18711 29348 18767 29404
rect 18767 29348 18771 29404
rect 18707 29344 18771 29348
rect 18787 29404 18851 29408
rect 18787 29348 18791 29404
rect 18791 29348 18847 29404
rect 18847 29348 18851 29404
rect 18787 29344 18851 29348
rect 18867 29404 18931 29408
rect 18867 29348 18871 29404
rect 18871 29348 18927 29404
rect 18927 29348 18931 29404
rect 18867 29344 18931 29348
rect 18947 29404 19011 29408
rect 18947 29348 18951 29404
rect 18951 29348 19007 29404
rect 19007 29348 19011 29404
rect 18947 29344 19011 29348
rect 3171 28860 3235 28864
rect 3171 28804 3175 28860
rect 3175 28804 3231 28860
rect 3231 28804 3235 28860
rect 3171 28800 3235 28804
rect 3251 28860 3315 28864
rect 3251 28804 3255 28860
rect 3255 28804 3311 28860
rect 3311 28804 3315 28860
rect 3251 28800 3315 28804
rect 3331 28860 3395 28864
rect 3331 28804 3335 28860
rect 3335 28804 3391 28860
rect 3391 28804 3395 28860
rect 3331 28800 3395 28804
rect 3411 28860 3475 28864
rect 3411 28804 3415 28860
rect 3415 28804 3471 28860
rect 3471 28804 3475 28860
rect 3411 28800 3475 28804
rect 7610 28860 7674 28864
rect 7610 28804 7614 28860
rect 7614 28804 7670 28860
rect 7670 28804 7674 28860
rect 7610 28800 7674 28804
rect 7690 28860 7754 28864
rect 7690 28804 7694 28860
rect 7694 28804 7750 28860
rect 7750 28804 7754 28860
rect 7690 28800 7754 28804
rect 7770 28860 7834 28864
rect 7770 28804 7774 28860
rect 7774 28804 7830 28860
rect 7830 28804 7834 28860
rect 7770 28800 7834 28804
rect 7850 28860 7914 28864
rect 7850 28804 7854 28860
rect 7854 28804 7910 28860
rect 7910 28804 7914 28860
rect 7850 28800 7914 28804
rect 12049 28860 12113 28864
rect 12049 28804 12053 28860
rect 12053 28804 12109 28860
rect 12109 28804 12113 28860
rect 12049 28800 12113 28804
rect 12129 28860 12193 28864
rect 12129 28804 12133 28860
rect 12133 28804 12189 28860
rect 12189 28804 12193 28860
rect 12129 28800 12193 28804
rect 12209 28860 12273 28864
rect 12209 28804 12213 28860
rect 12213 28804 12269 28860
rect 12269 28804 12273 28860
rect 12209 28800 12273 28804
rect 12289 28860 12353 28864
rect 12289 28804 12293 28860
rect 12293 28804 12349 28860
rect 12349 28804 12353 28860
rect 12289 28800 12353 28804
rect 16488 28860 16552 28864
rect 16488 28804 16492 28860
rect 16492 28804 16548 28860
rect 16548 28804 16552 28860
rect 16488 28800 16552 28804
rect 16568 28860 16632 28864
rect 16568 28804 16572 28860
rect 16572 28804 16628 28860
rect 16628 28804 16632 28860
rect 16568 28800 16632 28804
rect 16648 28860 16712 28864
rect 16648 28804 16652 28860
rect 16652 28804 16708 28860
rect 16708 28804 16712 28860
rect 16648 28800 16712 28804
rect 16728 28860 16792 28864
rect 16728 28804 16732 28860
rect 16732 28804 16788 28860
rect 16788 28804 16792 28860
rect 16728 28800 16792 28804
rect 5390 28316 5454 28320
rect 5390 28260 5394 28316
rect 5394 28260 5450 28316
rect 5450 28260 5454 28316
rect 5390 28256 5454 28260
rect 5470 28316 5534 28320
rect 5470 28260 5474 28316
rect 5474 28260 5530 28316
rect 5530 28260 5534 28316
rect 5470 28256 5534 28260
rect 5550 28316 5614 28320
rect 5550 28260 5554 28316
rect 5554 28260 5610 28316
rect 5610 28260 5614 28316
rect 5550 28256 5614 28260
rect 5630 28316 5694 28320
rect 5630 28260 5634 28316
rect 5634 28260 5690 28316
rect 5690 28260 5694 28316
rect 5630 28256 5694 28260
rect 9829 28316 9893 28320
rect 9829 28260 9833 28316
rect 9833 28260 9889 28316
rect 9889 28260 9893 28316
rect 9829 28256 9893 28260
rect 9909 28316 9973 28320
rect 9909 28260 9913 28316
rect 9913 28260 9969 28316
rect 9969 28260 9973 28316
rect 9909 28256 9973 28260
rect 9989 28316 10053 28320
rect 9989 28260 9993 28316
rect 9993 28260 10049 28316
rect 10049 28260 10053 28316
rect 9989 28256 10053 28260
rect 10069 28316 10133 28320
rect 10069 28260 10073 28316
rect 10073 28260 10129 28316
rect 10129 28260 10133 28316
rect 10069 28256 10133 28260
rect 14268 28316 14332 28320
rect 14268 28260 14272 28316
rect 14272 28260 14328 28316
rect 14328 28260 14332 28316
rect 14268 28256 14332 28260
rect 14348 28316 14412 28320
rect 14348 28260 14352 28316
rect 14352 28260 14408 28316
rect 14408 28260 14412 28316
rect 14348 28256 14412 28260
rect 14428 28316 14492 28320
rect 14428 28260 14432 28316
rect 14432 28260 14488 28316
rect 14488 28260 14492 28316
rect 14428 28256 14492 28260
rect 14508 28316 14572 28320
rect 14508 28260 14512 28316
rect 14512 28260 14568 28316
rect 14568 28260 14572 28316
rect 14508 28256 14572 28260
rect 18707 28316 18771 28320
rect 18707 28260 18711 28316
rect 18711 28260 18767 28316
rect 18767 28260 18771 28316
rect 18707 28256 18771 28260
rect 18787 28316 18851 28320
rect 18787 28260 18791 28316
rect 18791 28260 18847 28316
rect 18847 28260 18851 28316
rect 18787 28256 18851 28260
rect 18867 28316 18931 28320
rect 18867 28260 18871 28316
rect 18871 28260 18927 28316
rect 18927 28260 18931 28316
rect 18867 28256 18931 28260
rect 18947 28316 19011 28320
rect 18947 28260 18951 28316
rect 18951 28260 19007 28316
rect 19007 28260 19011 28316
rect 18947 28256 19011 28260
rect 3171 27772 3235 27776
rect 3171 27716 3175 27772
rect 3175 27716 3231 27772
rect 3231 27716 3235 27772
rect 3171 27712 3235 27716
rect 3251 27772 3315 27776
rect 3251 27716 3255 27772
rect 3255 27716 3311 27772
rect 3311 27716 3315 27772
rect 3251 27712 3315 27716
rect 3331 27772 3395 27776
rect 3331 27716 3335 27772
rect 3335 27716 3391 27772
rect 3391 27716 3395 27772
rect 3331 27712 3395 27716
rect 3411 27772 3475 27776
rect 3411 27716 3415 27772
rect 3415 27716 3471 27772
rect 3471 27716 3475 27772
rect 3411 27712 3475 27716
rect 7610 27772 7674 27776
rect 7610 27716 7614 27772
rect 7614 27716 7670 27772
rect 7670 27716 7674 27772
rect 7610 27712 7674 27716
rect 7690 27772 7754 27776
rect 7690 27716 7694 27772
rect 7694 27716 7750 27772
rect 7750 27716 7754 27772
rect 7690 27712 7754 27716
rect 7770 27772 7834 27776
rect 7770 27716 7774 27772
rect 7774 27716 7830 27772
rect 7830 27716 7834 27772
rect 7770 27712 7834 27716
rect 7850 27772 7914 27776
rect 7850 27716 7854 27772
rect 7854 27716 7910 27772
rect 7910 27716 7914 27772
rect 7850 27712 7914 27716
rect 12049 27772 12113 27776
rect 12049 27716 12053 27772
rect 12053 27716 12109 27772
rect 12109 27716 12113 27772
rect 12049 27712 12113 27716
rect 12129 27772 12193 27776
rect 12129 27716 12133 27772
rect 12133 27716 12189 27772
rect 12189 27716 12193 27772
rect 12129 27712 12193 27716
rect 12209 27772 12273 27776
rect 12209 27716 12213 27772
rect 12213 27716 12269 27772
rect 12269 27716 12273 27772
rect 12209 27712 12273 27716
rect 12289 27772 12353 27776
rect 12289 27716 12293 27772
rect 12293 27716 12349 27772
rect 12349 27716 12353 27772
rect 12289 27712 12353 27716
rect 16488 27772 16552 27776
rect 16488 27716 16492 27772
rect 16492 27716 16548 27772
rect 16548 27716 16552 27772
rect 16488 27712 16552 27716
rect 16568 27772 16632 27776
rect 16568 27716 16572 27772
rect 16572 27716 16628 27772
rect 16628 27716 16632 27772
rect 16568 27712 16632 27716
rect 16648 27772 16712 27776
rect 16648 27716 16652 27772
rect 16652 27716 16708 27772
rect 16708 27716 16712 27772
rect 16648 27712 16712 27716
rect 16728 27772 16792 27776
rect 16728 27716 16732 27772
rect 16732 27716 16788 27772
rect 16788 27716 16792 27772
rect 16728 27712 16792 27716
rect 5390 27228 5454 27232
rect 5390 27172 5394 27228
rect 5394 27172 5450 27228
rect 5450 27172 5454 27228
rect 5390 27168 5454 27172
rect 5470 27228 5534 27232
rect 5470 27172 5474 27228
rect 5474 27172 5530 27228
rect 5530 27172 5534 27228
rect 5470 27168 5534 27172
rect 5550 27228 5614 27232
rect 5550 27172 5554 27228
rect 5554 27172 5610 27228
rect 5610 27172 5614 27228
rect 5550 27168 5614 27172
rect 5630 27228 5694 27232
rect 5630 27172 5634 27228
rect 5634 27172 5690 27228
rect 5690 27172 5694 27228
rect 5630 27168 5694 27172
rect 9829 27228 9893 27232
rect 9829 27172 9833 27228
rect 9833 27172 9889 27228
rect 9889 27172 9893 27228
rect 9829 27168 9893 27172
rect 9909 27228 9973 27232
rect 9909 27172 9913 27228
rect 9913 27172 9969 27228
rect 9969 27172 9973 27228
rect 9909 27168 9973 27172
rect 9989 27228 10053 27232
rect 9989 27172 9993 27228
rect 9993 27172 10049 27228
rect 10049 27172 10053 27228
rect 9989 27168 10053 27172
rect 10069 27228 10133 27232
rect 10069 27172 10073 27228
rect 10073 27172 10129 27228
rect 10129 27172 10133 27228
rect 10069 27168 10133 27172
rect 14268 27228 14332 27232
rect 14268 27172 14272 27228
rect 14272 27172 14328 27228
rect 14328 27172 14332 27228
rect 14268 27168 14332 27172
rect 14348 27228 14412 27232
rect 14348 27172 14352 27228
rect 14352 27172 14408 27228
rect 14408 27172 14412 27228
rect 14348 27168 14412 27172
rect 14428 27228 14492 27232
rect 14428 27172 14432 27228
rect 14432 27172 14488 27228
rect 14488 27172 14492 27228
rect 14428 27168 14492 27172
rect 14508 27228 14572 27232
rect 14508 27172 14512 27228
rect 14512 27172 14568 27228
rect 14568 27172 14572 27228
rect 14508 27168 14572 27172
rect 18707 27228 18771 27232
rect 18707 27172 18711 27228
rect 18711 27172 18767 27228
rect 18767 27172 18771 27228
rect 18707 27168 18771 27172
rect 18787 27228 18851 27232
rect 18787 27172 18791 27228
rect 18791 27172 18847 27228
rect 18847 27172 18851 27228
rect 18787 27168 18851 27172
rect 18867 27228 18931 27232
rect 18867 27172 18871 27228
rect 18871 27172 18927 27228
rect 18927 27172 18931 27228
rect 18867 27168 18931 27172
rect 18947 27228 19011 27232
rect 18947 27172 18951 27228
rect 18951 27172 19007 27228
rect 19007 27172 19011 27228
rect 18947 27168 19011 27172
rect 3171 26684 3235 26688
rect 3171 26628 3175 26684
rect 3175 26628 3231 26684
rect 3231 26628 3235 26684
rect 3171 26624 3235 26628
rect 3251 26684 3315 26688
rect 3251 26628 3255 26684
rect 3255 26628 3311 26684
rect 3311 26628 3315 26684
rect 3251 26624 3315 26628
rect 3331 26684 3395 26688
rect 3331 26628 3335 26684
rect 3335 26628 3391 26684
rect 3391 26628 3395 26684
rect 3331 26624 3395 26628
rect 3411 26684 3475 26688
rect 3411 26628 3415 26684
rect 3415 26628 3471 26684
rect 3471 26628 3475 26684
rect 3411 26624 3475 26628
rect 7610 26684 7674 26688
rect 7610 26628 7614 26684
rect 7614 26628 7670 26684
rect 7670 26628 7674 26684
rect 7610 26624 7674 26628
rect 7690 26684 7754 26688
rect 7690 26628 7694 26684
rect 7694 26628 7750 26684
rect 7750 26628 7754 26684
rect 7690 26624 7754 26628
rect 7770 26684 7834 26688
rect 7770 26628 7774 26684
rect 7774 26628 7830 26684
rect 7830 26628 7834 26684
rect 7770 26624 7834 26628
rect 7850 26684 7914 26688
rect 7850 26628 7854 26684
rect 7854 26628 7910 26684
rect 7910 26628 7914 26684
rect 7850 26624 7914 26628
rect 12049 26684 12113 26688
rect 12049 26628 12053 26684
rect 12053 26628 12109 26684
rect 12109 26628 12113 26684
rect 12049 26624 12113 26628
rect 12129 26684 12193 26688
rect 12129 26628 12133 26684
rect 12133 26628 12189 26684
rect 12189 26628 12193 26684
rect 12129 26624 12193 26628
rect 12209 26684 12273 26688
rect 12209 26628 12213 26684
rect 12213 26628 12269 26684
rect 12269 26628 12273 26684
rect 12209 26624 12273 26628
rect 12289 26684 12353 26688
rect 12289 26628 12293 26684
rect 12293 26628 12349 26684
rect 12349 26628 12353 26684
rect 12289 26624 12353 26628
rect 16488 26684 16552 26688
rect 16488 26628 16492 26684
rect 16492 26628 16548 26684
rect 16548 26628 16552 26684
rect 16488 26624 16552 26628
rect 16568 26684 16632 26688
rect 16568 26628 16572 26684
rect 16572 26628 16628 26684
rect 16628 26628 16632 26684
rect 16568 26624 16632 26628
rect 16648 26684 16712 26688
rect 16648 26628 16652 26684
rect 16652 26628 16708 26684
rect 16708 26628 16712 26684
rect 16648 26624 16712 26628
rect 16728 26684 16792 26688
rect 16728 26628 16732 26684
rect 16732 26628 16788 26684
rect 16788 26628 16792 26684
rect 16728 26624 16792 26628
rect 5390 26140 5454 26144
rect 5390 26084 5394 26140
rect 5394 26084 5450 26140
rect 5450 26084 5454 26140
rect 5390 26080 5454 26084
rect 5470 26140 5534 26144
rect 5470 26084 5474 26140
rect 5474 26084 5530 26140
rect 5530 26084 5534 26140
rect 5470 26080 5534 26084
rect 5550 26140 5614 26144
rect 5550 26084 5554 26140
rect 5554 26084 5610 26140
rect 5610 26084 5614 26140
rect 5550 26080 5614 26084
rect 5630 26140 5694 26144
rect 5630 26084 5634 26140
rect 5634 26084 5690 26140
rect 5690 26084 5694 26140
rect 5630 26080 5694 26084
rect 9829 26140 9893 26144
rect 9829 26084 9833 26140
rect 9833 26084 9889 26140
rect 9889 26084 9893 26140
rect 9829 26080 9893 26084
rect 9909 26140 9973 26144
rect 9909 26084 9913 26140
rect 9913 26084 9969 26140
rect 9969 26084 9973 26140
rect 9909 26080 9973 26084
rect 9989 26140 10053 26144
rect 9989 26084 9993 26140
rect 9993 26084 10049 26140
rect 10049 26084 10053 26140
rect 9989 26080 10053 26084
rect 10069 26140 10133 26144
rect 10069 26084 10073 26140
rect 10073 26084 10129 26140
rect 10129 26084 10133 26140
rect 10069 26080 10133 26084
rect 14268 26140 14332 26144
rect 14268 26084 14272 26140
rect 14272 26084 14328 26140
rect 14328 26084 14332 26140
rect 14268 26080 14332 26084
rect 14348 26140 14412 26144
rect 14348 26084 14352 26140
rect 14352 26084 14408 26140
rect 14408 26084 14412 26140
rect 14348 26080 14412 26084
rect 14428 26140 14492 26144
rect 14428 26084 14432 26140
rect 14432 26084 14488 26140
rect 14488 26084 14492 26140
rect 14428 26080 14492 26084
rect 14508 26140 14572 26144
rect 14508 26084 14512 26140
rect 14512 26084 14568 26140
rect 14568 26084 14572 26140
rect 14508 26080 14572 26084
rect 18707 26140 18771 26144
rect 18707 26084 18711 26140
rect 18711 26084 18767 26140
rect 18767 26084 18771 26140
rect 18707 26080 18771 26084
rect 18787 26140 18851 26144
rect 18787 26084 18791 26140
rect 18791 26084 18847 26140
rect 18847 26084 18851 26140
rect 18787 26080 18851 26084
rect 18867 26140 18931 26144
rect 18867 26084 18871 26140
rect 18871 26084 18927 26140
rect 18927 26084 18931 26140
rect 18867 26080 18931 26084
rect 18947 26140 19011 26144
rect 18947 26084 18951 26140
rect 18951 26084 19007 26140
rect 19007 26084 19011 26140
rect 18947 26080 19011 26084
rect 3171 25596 3235 25600
rect 3171 25540 3175 25596
rect 3175 25540 3231 25596
rect 3231 25540 3235 25596
rect 3171 25536 3235 25540
rect 3251 25596 3315 25600
rect 3251 25540 3255 25596
rect 3255 25540 3311 25596
rect 3311 25540 3315 25596
rect 3251 25536 3315 25540
rect 3331 25596 3395 25600
rect 3331 25540 3335 25596
rect 3335 25540 3391 25596
rect 3391 25540 3395 25596
rect 3331 25536 3395 25540
rect 3411 25596 3475 25600
rect 3411 25540 3415 25596
rect 3415 25540 3471 25596
rect 3471 25540 3475 25596
rect 3411 25536 3475 25540
rect 7610 25596 7674 25600
rect 7610 25540 7614 25596
rect 7614 25540 7670 25596
rect 7670 25540 7674 25596
rect 7610 25536 7674 25540
rect 7690 25596 7754 25600
rect 7690 25540 7694 25596
rect 7694 25540 7750 25596
rect 7750 25540 7754 25596
rect 7690 25536 7754 25540
rect 7770 25596 7834 25600
rect 7770 25540 7774 25596
rect 7774 25540 7830 25596
rect 7830 25540 7834 25596
rect 7770 25536 7834 25540
rect 7850 25596 7914 25600
rect 7850 25540 7854 25596
rect 7854 25540 7910 25596
rect 7910 25540 7914 25596
rect 7850 25536 7914 25540
rect 12049 25596 12113 25600
rect 12049 25540 12053 25596
rect 12053 25540 12109 25596
rect 12109 25540 12113 25596
rect 12049 25536 12113 25540
rect 12129 25596 12193 25600
rect 12129 25540 12133 25596
rect 12133 25540 12189 25596
rect 12189 25540 12193 25596
rect 12129 25536 12193 25540
rect 12209 25596 12273 25600
rect 12209 25540 12213 25596
rect 12213 25540 12269 25596
rect 12269 25540 12273 25596
rect 12209 25536 12273 25540
rect 12289 25596 12353 25600
rect 12289 25540 12293 25596
rect 12293 25540 12349 25596
rect 12349 25540 12353 25596
rect 12289 25536 12353 25540
rect 16488 25596 16552 25600
rect 16488 25540 16492 25596
rect 16492 25540 16548 25596
rect 16548 25540 16552 25596
rect 16488 25536 16552 25540
rect 16568 25596 16632 25600
rect 16568 25540 16572 25596
rect 16572 25540 16628 25596
rect 16628 25540 16632 25596
rect 16568 25536 16632 25540
rect 16648 25596 16712 25600
rect 16648 25540 16652 25596
rect 16652 25540 16708 25596
rect 16708 25540 16712 25596
rect 16648 25536 16712 25540
rect 16728 25596 16792 25600
rect 16728 25540 16732 25596
rect 16732 25540 16788 25596
rect 16788 25540 16792 25596
rect 16728 25536 16792 25540
rect 5390 25052 5454 25056
rect 5390 24996 5394 25052
rect 5394 24996 5450 25052
rect 5450 24996 5454 25052
rect 5390 24992 5454 24996
rect 5470 25052 5534 25056
rect 5470 24996 5474 25052
rect 5474 24996 5530 25052
rect 5530 24996 5534 25052
rect 5470 24992 5534 24996
rect 5550 25052 5614 25056
rect 5550 24996 5554 25052
rect 5554 24996 5610 25052
rect 5610 24996 5614 25052
rect 5550 24992 5614 24996
rect 5630 25052 5694 25056
rect 5630 24996 5634 25052
rect 5634 24996 5690 25052
rect 5690 24996 5694 25052
rect 5630 24992 5694 24996
rect 9829 25052 9893 25056
rect 9829 24996 9833 25052
rect 9833 24996 9889 25052
rect 9889 24996 9893 25052
rect 9829 24992 9893 24996
rect 9909 25052 9973 25056
rect 9909 24996 9913 25052
rect 9913 24996 9969 25052
rect 9969 24996 9973 25052
rect 9909 24992 9973 24996
rect 9989 25052 10053 25056
rect 9989 24996 9993 25052
rect 9993 24996 10049 25052
rect 10049 24996 10053 25052
rect 9989 24992 10053 24996
rect 10069 25052 10133 25056
rect 10069 24996 10073 25052
rect 10073 24996 10129 25052
rect 10129 24996 10133 25052
rect 10069 24992 10133 24996
rect 14268 25052 14332 25056
rect 14268 24996 14272 25052
rect 14272 24996 14328 25052
rect 14328 24996 14332 25052
rect 14268 24992 14332 24996
rect 14348 25052 14412 25056
rect 14348 24996 14352 25052
rect 14352 24996 14408 25052
rect 14408 24996 14412 25052
rect 14348 24992 14412 24996
rect 14428 25052 14492 25056
rect 14428 24996 14432 25052
rect 14432 24996 14488 25052
rect 14488 24996 14492 25052
rect 14428 24992 14492 24996
rect 14508 25052 14572 25056
rect 14508 24996 14512 25052
rect 14512 24996 14568 25052
rect 14568 24996 14572 25052
rect 14508 24992 14572 24996
rect 18707 25052 18771 25056
rect 18707 24996 18711 25052
rect 18711 24996 18767 25052
rect 18767 24996 18771 25052
rect 18707 24992 18771 24996
rect 18787 25052 18851 25056
rect 18787 24996 18791 25052
rect 18791 24996 18847 25052
rect 18847 24996 18851 25052
rect 18787 24992 18851 24996
rect 18867 25052 18931 25056
rect 18867 24996 18871 25052
rect 18871 24996 18927 25052
rect 18927 24996 18931 25052
rect 18867 24992 18931 24996
rect 18947 25052 19011 25056
rect 18947 24996 18951 25052
rect 18951 24996 19007 25052
rect 19007 24996 19011 25052
rect 18947 24992 19011 24996
rect 3171 24508 3235 24512
rect 3171 24452 3175 24508
rect 3175 24452 3231 24508
rect 3231 24452 3235 24508
rect 3171 24448 3235 24452
rect 3251 24508 3315 24512
rect 3251 24452 3255 24508
rect 3255 24452 3311 24508
rect 3311 24452 3315 24508
rect 3251 24448 3315 24452
rect 3331 24508 3395 24512
rect 3331 24452 3335 24508
rect 3335 24452 3391 24508
rect 3391 24452 3395 24508
rect 3331 24448 3395 24452
rect 3411 24508 3475 24512
rect 3411 24452 3415 24508
rect 3415 24452 3471 24508
rect 3471 24452 3475 24508
rect 3411 24448 3475 24452
rect 7610 24508 7674 24512
rect 7610 24452 7614 24508
rect 7614 24452 7670 24508
rect 7670 24452 7674 24508
rect 7610 24448 7674 24452
rect 7690 24508 7754 24512
rect 7690 24452 7694 24508
rect 7694 24452 7750 24508
rect 7750 24452 7754 24508
rect 7690 24448 7754 24452
rect 7770 24508 7834 24512
rect 7770 24452 7774 24508
rect 7774 24452 7830 24508
rect 7830 24452 7834 24508
rect 7770 24448 7834 24452
rect 7850 24508 7914 24512
rect 7850 24452 7854 24508
rect 7854 24452 7910 24508
rect 7910 24452 7914 24508
rect 7850 24448 7914 24452
rect 12049 24508 12113 24512
rect 12049 24452 12053 24508
rect 12053 24452 12109 24508
rect 12109 24452 12113 24508
rect 12049 24448 12113 24452
rect 12129 24508 12193 24512
rect 12129 24452 12133 24508
rect 12133 24452 12189 24508
rect 12189 24452 12193 24508
rect 12129 24448 12193 24452
rect 12209 24508 12273 24512
rect 12209 24452 12213 24508
rect 12213 24452 12269 24508
rect 12269 24452 12273 24508
rect 12209 24448 12273 24452
rect 12289 24508 12353 24512
rect 12289 24452 12293 24508
rect 12293 24452 12349 24508
rect 12349 24452 12353 24508
rect 12289 24448 12353 24452
rect 16488 24508 16552 24512
rect 16488 24452 16492 24508
rect 16492 24452 16548 24508
rect 16548 24452 16552 24508
rect 16488 24448 16552 24452
rect 16568 24508 16632 24512
rect 16568 24452 16572 24508
rect 16572 24452 16628 24508
rect 16628 24452 16632 24508
rect 16568 24448 16632 24452
rect 16648 24508 16712 24512
rect 16648 24452 16652 24508
rect 16652 24452 16708 24508
rect 16708 24452 16712 24508
rect 16648 24448 16712 24452
rect 16728 24508 16792 24512
rect 16728 24452 16732 24508
rect 16732 24452 16788 24508
rect 16788 24452 16792 24508
rect 16728 24448 16792 24452
rect 5390 23964 5454 23968
rect 5390 23908 5394 23964
rect 5394 23908 5450 23964
rect 5450 23908 5454 23964
rect 5390 23904 5454 23908
rect 5470 23964 5534 23968
rect 5470 23908 5474 23964
rect 5474 23908 5530 23964
rect 5530 23908 5534 23964
rect 5470 23904 5534 23908
rect 5550 23964 5614 23968
rect 5550 23908 5554 23964
rect 5554 23908 5610 23964
rect 5610 23908 5614 23964
rect 5550 23904 5614 23908
rect 5630 23964 5694 23968
rect 5630 23908 5634 23964
rect 5634 23908 5690 23964
rect 5690 23908 5694 23964
rect 5630 23904 5694 23908
rect 9829 23964 9893 23968
rect 9829 23908 9833 23964
rect 9833 23908 9889 23964
rect 9889 23908 9893 23964
rect 9829 23904 9893 23908
rect 9909 23964 9973 23968
rect 9909 23908 9913 23964
rect 9913 23908 9969 23964
rect 9969 23908 9973 23964
rect 9909 23904 9973 23908
rect 9989 23964 10053 23968
rect 9989 23908 9993 23964
rect 9993 23908 10049 23964
rect 10049 23908 10053 23964
rect 9989 23904 10053 23908
rect 10069 23964 10133 23968
rect 10069 23908 10073 23964
rect 10073 23908 10129 23964
rect 10129 23908 10133 23964
rect 10069 23904 10133 23908
rect 14268 23964 14332 23968
rect 14268 23908 14272 23964
rect 14272 23908 14328 23964
rect 14328 23908 14332 23964
rect 14268 23904 14332 23908
rect 14348 23964 14412 23968
rect 14348 23908 14352 23964
rect 14352 23908 14408 23964
rect 14408 23908 14412 23964
rect 14348 23904 14412 23908
rect 14428 23964 14492 23968
rect 14428 23908 14432 23964
rect 14432 23908 14488 23964
rect 14488 23908 14492 23964
rect 14428 23904 14492 23908
rect 14508 23964 14572 23968
rect 14508 23908 14512 23964
rect 14512 23908 14568 23964
rect 14568 23908 14572 23964
rect 14508 23904 14572 23908
rect 18707 23964 18771 23968
rect 18707 23908 18711 23964
rect 18711 23908 18767 23964
rect 18767 23908 18771 23964
rect 18707 23904 18771 23908
rect 18787 23964 18851 23968
rect 18787 23908 18791 23964
rect 18791 23908 18847 23964
rect 18847 23908 18851 23964
rect 18787 23904 18851 23908
rect 18867 23964 18931 23968
rect 18867 23908 18871 23964
rect 18871 23908 18927 23964
rect 18927 23908 18931 23964
rect 18867 23904 18931 23908
rect 18947 23964 19011 23968
rect 18947 23908 18951 23964
rect 18951 23908 19007 23964
rect 19007 23908 19011 23964
rect 18947 23904 19011 23908
rect 3171 23420 3235 23424
rect 3171 23364 3175 23420
rect 3175 23364 3231 23420
rect 3231 23364 3235 23420
rect 3171 23360 3235 23364
rect 3251 23420 3315 23424
rect 3251 23364 3255 23420
rect 3255 23364 3311 23420
rect 3311 23364 3315 23420
rect 3251 23360 3315 23364
rect 3331 23420 3395 23424
rect 3331 23364 3335 23420
rect 3335 23364 3391 23420
rect 3391 23364 3395 23420
rect 3331 23360 3395 23364
rect 3411 23420 3475 23424
rect 3411 23364 3415 23420
rect 3415 23364 3471 23420
rect 3471 23364 3475 23420
rect 3411 23360 3475 23364
rect 7610 23420 7674 23424
rect 7610 23364 7614 23420
rect 7614 23364 7670 23420
rect 7670 23364 7674 23420
rect 7610 23360 7674 23364
rect 7690 23420 7754 23424
rect 7690 23364 7694 23420
rect 7694 23364 7750 23420
rect 7750 23364 7754 23420
rect 7690 23360 7754 23364
rect 7770 23420 7834 23424
rect 7770 23364 7774 23420
rect 7774 23364 7830 23420
rect 7830 23364 7834 23420
rect 7770 23360 7834 23364
rect 7850 23420 7914 23424
rect 7850 23364 7854 23420
rect 7854 23364 7910 23420
rect 7910 23364 7914 23420
rect 7850 23360 7914 23364
rect 12049 23420 12113 23424
rect 12049 23364 12053 23420
rect 12053 23364 12109 23420
rect 12109 23364 12113 23420
rect 12049 23360 12113 23364
rect 12129 23420 12193 23424
rect 12129 23364 12133 23420
rect 12133 23364 12189 23420
rect 12189 23364 12193 23420
rect 12129 23360 12193 23364
rect 12209 23420 12273 23424
rect 12209 23364 12213 23420
rect 12213 23364 12269 23420
rect 12269 23364 12273 23420
rect 12209 23360 12273 23364
rect 12289 23420 12353 23424
rect 12289 23364 12293 23420
rect 12293 23364 12349 23420
rect 12349 23364 12353 23420
rect 12289 23360 12353 23364
rect 16488 23420 16552 23424
rect 16488 23364 16492 23420
rect 16492 23364 16548 23420
rect 16548 23364 16552 23420
rect 16488 23360 16552 23364
rect 16568 23420 16632 23424
rect 16568 23364 16572 23420
rect 16572 23364 16628 23420
rect 16628 23364 16632 23420
rect 16568 23360 16632 23364
rect 16648 23420 16712 23424
rect 16648 23364 16652 23420
rect 16652 23364 16708 23420
rect 16708 23364 16712 23420
rect 16648 23360 16712 23364
rect 16728 23420 16792 23424
rect 16728 23364 16732 23420
rect 16732 23364 16788 23420
rect 16788 23364 16792 23420
rect 16728 23360 16792 23364
rect 5390 22876 5454 22880
rect 5390 22820 5394 22876
rect 5394 22820 5450 22876
rect 5450 22820 5454 22876
rect 5390 22816 5454 22820
rect 5470 22876 5534 22880
rect 5470 22820 5474 22876
rect 5474 22820 5530 22876
rect 5530 22820 5534 22876
rect 5470 22816 5534 22820
rect 5550 22876 5614 22880
rect 5550 22820 5554 22876
rect 5554 22820 5610 22876
rect 5610 22820 5614 22876
rect 5550 22816 5614 22820
rect 5630 22876 5694 22880
rect 5630 22820 5634 22876
rect 5634 22820 5690 22876
rect 5690 22820 5694 22876
rect 5630 22816 5694 22820
rect 9829 22876 9893 22880
rect 9829 22820 9833 22876
rect 9833 22820 9889 22876
rect 9889 22820 9893 22876
rect 9829 22816 9893 22820
rect 9909 22876 9973 22880
rect 9909 22820 9913 22876
rect 9913 22820 9969 22876
rect 9969 22820 9973 22876
rect 9909 22816 9973 22820
rect 9989 22876 10053 22880
rect 9989 22820 9993 22876
rect 9993 22820 10049 22876
rect 10049 22820 10053 22876
rect 9989 22816 10053 22820
rect 10069 22876 10133 22880
rect 10069 22820 10073 22876
rect 10073 22820 10129 22876
rect 10129 22820 10133 22876
rect 10069 22816 10133 22820
rect 14268 22876 14332 22880
rect 14268 22820 14272 22876
rect 14272 22820 14328 22876
rect 14328 22820 14332 22876
rect 14268 22816 14332 22820
rect 14348 22876 14412 22880
rect 14348 22820 14352 22876
rect 14352 22820 14408 22876
rect 14408 22820 14412 22876
rect 14348 22816 14412 22820
rect 14428 22876 14492 22880
rect 14428 22820 14432 22876
rect 14432 22820 14488 22876
rect 14488 22820 14492 22876
rect 14428 22816 14492 22820
rect 14508 22876 14572 22880
rect 14508 22820 14512 22876
rect 14512 22820 14568 22876
rect 14568 22820 14572 22876
rect 14508 22816 14572 22820
rect 18707 22876 18771 22880
rect 18707 22820 18711 22876
rect 18711 22820 18767 22876
rect 18767 22820 18771 22876
rect 18707 22816 18771 22820
rect 18787 22876 18851 22880
rect 18787 22820 18791 22876
rect 18791 22820 18847 22876
rect 18847 22820 18851 22876
rect 18787 22816 18851 22820
rect 18867 22876 18931 22880
rect 18867 22820 18871 22876
rect 18871 22820 18927 22876
rect 18927 22820 18931 22876
rect 18867 22816 18931 22820
rect 18947 22876 19011 22880
rect 18947 22820 18951 22876
rect 18951 22820 19007 22876
rect 19007 22820 19011 22876
rect 18947 22816 19011 22820
rect 3171 22332 3235 22336
rect 3171 22276 3175 22332
rect 3175 22276 3231 22332
rect 3231 22276 3235 22332
rect 3171 22272 3235 22276
rect 3251 22332 3315 22336
rect 3251 22276 3255 22332
rect 3255 22276 3311 22332
rect 3311 22276 3315 22332
rect 3251 22272 3315 22276
rect 3331 22332 3395 22336
rect 3331 22276 3335 22332
rect 3335 22276 3391 22332
rect 3391 22276 3395 22332
rect 3331 22272 3395 22276
rect 3411 22332 3475 22336
rect 3411 22276 3415 22332
rect 3415 22276 3471 22332
rect 3471 22276 3475 22332
rect 3411 22272 3475 22276
rect 7610 22332 7674 22336
rect 7610 22276 7614 22332
rect 7614 22276 7670 22332
rect 7670 22276 7674 22332
rect 7610 22272 7674 22276
rect 7690 22332 7754 22336
rect 7690 22276 7694 22332
rect 7694 22276 7750 22332
rect 7750 22276 7754 22332
rect 7690 22272 7754 22276
rect 7770 22332 7834 22336
rect 7770 22276 7774 22332
rect 7774 22276 7830 22332
rect 7830 22276 7834 22332
rect 7770 22272 7834 22276
rect 7850 22332 7914 22336
rect 7850 22276 7854 22332
rect 7854 22276 7910 22332
rect 7910 22276 7914 22332
rect 7850 22272 7914 22276
rect 12049 22332 12113 22336
rect 12049 22276 12053 22332
rect 12053 22276 12109 22332
rect 12109 22276 12113 22332
rect 12049 22272 12113 22276
rect 12129 22332 12193 22336
rect 12129 22276 12133 22332
rect 12133 22276 12189 22332
rect 12189 22276 12193 22332
rect 12129 22272 12193 22276
rect 12209 22332 12273 22336
rect 12209 22276 12213 22332
rect 12213 22276 12269 22332
rect 12269 22276 12273 22332
rect 12209 22272 12273 22276
rect 12289 22332 12353 22336
rect 12289 22276 12293 22332
rect 12293 22276 12349 22332
rect 12349 22276 12353 22332
rect 12289 22272 12353 22276
rect 16488 22332 16552 22336
rect 16488 22276 16492 22332
rect 16492 22276 16548 22332
rect 16548 22276 16552 22332
rect 16488 22272 16552 22276
rect 16568 22332 16632 22336
rect 16568 22276 16572 22332
rect 16572 22276 16628 22332
rect 16628 22276 16632 22332
rect 16568 22272 16632 22276
rect 16648 22332 16712 22336
rect 16648 22276 16652 22332
rect 16652 22276 16708 22332
rect 16708 22276 16712 22332
rect 16648 22272 16712 22276
rect 16728 22332 16792 22336
rect 16728 22276 16732 22332
rect 16732 22276 16788 22332
rect 16788 22276 16792 22332
rect 16728 22272 16792 22276
rect 5390 21788 5454 21792
rect 5390 21732 5394 21788
rect 5394 21732 5450 21788
rect 5450 21732 5454 21788
rect 5390 21728 5454 21732
rect 5470 21788 5534 21792
rect 5470 21732 5474 21788
rect 5474 21732 5530 21788
rect 5530 21732 5534 21788
rect 5470 21728 5534 21732
rect 5550 21788 5614 21792
rect 5550 21732 5554 21788
rect 5554 21732 5610 21788
rect 5610 21732 5614 21788
rect 5550 21728 5614 21732
rect 5630 21788 5694 21792
rect 5630 21732 5634 21788
rect 5634 21732 5690 21788
rect 5690 21732 5694 21788
rect 5630 21728 5694 21732
rect 9829 21788 9893 21792
rect 9829 21732 9833 21788
rect 9833 21732 9889 21788
rect 9889 21732 9893 21788
rect 9829 21728 9893 21732
rect 9909 21788 9973 21792
rect 9909 21732 9913 21788
rect 9913 21732 9969 21788
rect 9969 21732 9973 21788
rect 9909 21728 9973 21732
rect 9989 21788 10053 21792
rect 9989 21732 9993 21788
rect 9993 21732 10049 21788
rect 10049 21732 10053 21788
rect 9989 21728 10053 21732
rect 10069 21788 10133 21792
rect 10069 21732 10073 21788
rect 10073 21732 10129 21788
rect 10129 21732 10133 21788
rect 10069 21728 10133 21732
rect 14268 21788 14332 21792
rect 14268 21732 14272 21788
rect 14272 21732 14328 21788
rect 14328 21732 14332 21788
rect 14268 21728 14332 21732
rect 14348 21788 14412 21792
rect 14348 21732 14352 21788
rect 14352 21732 14408 21788
rect 14408 21732 14412 21788
rect 14348 21728 14412 21732
rect 14428 21788 14492 21792
rect 14428 21732 14432 21788
rect 14432 21732 14488 21788
rect 14488 21732 14492 21788
rect 14428 21728 14492 21732
rect 14508 21788 14572 21792
rect 14508 21732 14512 21788
rect 14512 21732 14568 21788
rect 14568 21732 14572 21788
rect 14508 21728 14572 21732
rect 18707 21788 18771 21792
rect 18707 21732 18711 21788
rect 18711 21732 18767 21788
rect 18767 21732 18771 21788
rect 18707 21728 18771 21732
rect 18787 21788 18851 21792
rect 18787 21732 18791 21788
rect 18791 21732 18847 21788
rect 18847 21732 18851 21788
rect 18787 21728 18851 21732
rect 18867 21788 18931 21792
rect 18867 21732 18871 21788
rect 18871 21732 18927 21788
rect 18927 21732 18931 21788
rect 18867 21728 18931 21732
rect 18947 21788 19011 21792
rect 18947 21732 18951 21788
rect 18951 21732 19007 21788
rect 19007 21732 19011 21788
rect 18947 21728 19011 21732
rect 3171 21244 3235 21248
rect 3171 21188 3175 21244
rect 3175 21188 3231 21244
rect 3231 21188 3235 21244
rect 3171 21184 3235 21188
rect 3251 21244 3315 21248
rect 3251 21188 3255 21244
rect 3255 21188 3311 21244
rect 3311 21188 3315 21244
rect 3251 21184 3315 21188
rect 3331 21244 3395 21248
rect 3331 21188 3335 21244
rect 3335 21188 3391 21244
rect 3391 21188 3395 21244
rect 3331 21184 3395 21188
rect 3411 21244 3475 21248
rect 3411 21188 3415 21244
rect 3415 21188 3471 21244
rect 3471 21188 3475 21244
rect 3411 21184 3475 21188
rect 7610 21244 7674 21248
rect 7610 21188 7614 21244
rect 7614 21188 7670 21244
rect 7670 21188 7674 21244
rect 7610 21184 7674 21188
rect 7690 21244 7754 21248
rect 7690 21188 7694 21244
rect 7694 21188 7750 21244
rect 7750 21188 7754 21244
rect 7690 21184 7754 21188
rect 7770 21244 7834 21248
rect 7770 21188 7774 21244
rect 7774 21188 7830 21244
rect 7830 21188 7834 21244
rect 7770 21184 7834 21188
rect 7850 21244 7914 21248
rect 7850 21188 7854 21244
rect 7854 21188 7910 21244
rect 7910 21188 7914 21244
rect 7850 21184 7914 21188
rect 12049 21244 12113 21248
rect 12049 21188 12053 21244
rect 12053 21188 12109 21244
rect 12109 21188 12113 21244
rect 12049 21184 12113 21188
rect 12129 21244 12193 21248
rect 12129 21188 12133 21244
rect 12133 21188 12189 21244
rect 12189 21188 12193 21244
rect 12129 21184 12193 21188
rect 12209 21244 12273 21248
rect 12209 21188 12213 21244
rect 12213 21188 12269 21244
rect 12269 21188 12273 21244
rect 12209 21184 12273 21188
rect 12289 21244 12353 21248
rect 12289 21188 12293 21244
rect 12293 21188 12349 21244
rect 12349 21188 12353 21244
rect 12289 21184 12353 21188
rect 16488 21244 16552 21248
rect 16488 21188 16492 21244
rect 16492 21188 16548 21244
rect 16548 21188 16552 21244
rect 16488 21184 16552 21188
rect 16568 21244 16632 21248
rect 16568 21188 16572 21244
rect 16572 21188 16628 21244
rect 16628 21188 16632 21244
rect 16568 21184 16632 21188
rect 16648 21244 16712 21248
rect 16648 21188 16652 21244
rect 16652 21188 16708 21244
rect 16708 21188 16712 21244
rect 16648 21184 16712 21188
rect 16728 21244 16792 21248
rect 16728 21188 16732 21244
rect 16732 21188 16788 21244
rect 16788 21188 16792 21244
rect 16728 21184 16792 21188
rect 5390 20700 5454 20704
rect 5390 20644 5394 20700
rect 5394 20644 5450 20700
rect 5450 20644 5454 20700
rect 5390 20640 5454 20644
rect 5470 20700 5534 20704
rect 5470 20644 5474 20700
rect 5474 20644 5530 20700
rect 5530 20644 5534 20700
rect 5470 20640 5534 20644
rect 5550 20700 5614 20704
rect 5550 20644 5554 20700
rect 5554 20644 5610 20700
rect 5610 20644 5614 20700
rect 5550 20640 5614 20644
rect 5630 20700 5694 20704
rect 5630 20644 5634 20700
rect 5634 20644 5690 20700
rect 5690 20644 5694 20700
rect 5630 20640 5694 20644
rect 9829 20700 9893 20704
rect 9829 20644 9833 20700
rect 9833 20644 9889 20700
rect 9889 20644 9893 20700
rect 9829 20640 9893 20644
rect 9909 20700 9973 20704
rect 9909 20644 9913 20700
rect 9913 20644 9969 20700
rect 9969 20644 9973 20700
rect 9909 20640 9973 20644
rect 9989 20700 10053 20704
rect 9989 20644 9993 20700
rect 9993 20644 10049 20700
rect 10049 20644 10053 20700
rect 9989 20640 10053 20644
rect 10069 20700 10133 20704
rect 10069 20644 10073 20700
rect 10073 20644 10129 20700
rect 10129 20644 10133 20700
rect 10069 20640 10133 20644
rect 14268 20700 14332 20704
rect 14268 20644 14272 20700
rect 14272 20644 14328 20700
rect 14328 20644 14332 20700
rect 14268 20640 14332 20644
rect 14348 20700 14412 20704
rect 14348 20644 14352 20700
rect 14352 20644 14408 20700
rect 14408 20644 14412 20700
rect 14348 20640 14412 20644
rect 14428 20700 14492 20704
rect 14428 20644 14432 20700
rect 14432 20644 14488 20700
rect 14488 20644 14492 20700
rect 14428 20640 14492 20644
rect 14508 20700 14572 20704
rect 14508 20644 14512 20700
rect 14512 20644 14568 20700
rect 14568 20644 14572 20700
rect 14508 20640 14572 20644
rect 18707 20700 18771 20704
rect 18707 20644 18711 20700
rect 18711 20644 18767 20700
rect 18767 20644 18771 20700
rect 18707 20640 18771 20644
rect 18787 20700 18851 20704
rect 18787 20644 18791 20700
rect 18791 20644 18847 20700
rect 18847 20644 18851 20700
rect 18787 20640 18851 20644
rect 18867 20700 18931 20704
rect 18867 20644 18871 20700
rect 18871 20644 18927 20700
rect 18927 20644 18931 20700
rect 18867 20640 18931 20644
rect 18947 20700 19011 20704
rect 18947 20644 18951 20700
rect 18951 20644 19007 20700
rect 19007 20644 19011 20700
rect 18947 20640 19011 20644
rect 3171 20156 3235 20160
rect 3171 20100 3175 20156
rect 3175 20100 3231 20156
rect 3231 20100 3235 20156
rect 3171 20096 3235 20100
rect 3251 20156 3315 20160
rect 3251 20100 3255 20156
rect 3255 20100 3311 20156
rect 3311 20100 3315 20156
rect 3251 20096 3315 20100
rect 3331 20156 3395 20160
rect 3331 20100 3335 20156
rect 3335 20100 3391 20156
rect 3391 20100 3395 20156
rect 3331 20096 3395 20100
rect 3411 20156 3475 20160
rect 3411 20100 3415 20156
rect 3415 20100 3471 20156
rect 3471 20100 3475 20156
rect 3411 20096 3475 20100
rect 7610 20156 7674 20160
rect 7610 20100 7614 20156
rect 7614 20100 7670 20156
rect 7670 20100 7674 20156
rect 7610 20096 7674 20100
rect 7690 20156 7754 20160
rect 7690 20100 7694 20156
rect 7694 20100 7750 20156
rect 7750 20100 7754 20156
rect 7690 20096 7754 20100
rect 7770 20156 7834 20160
rect 7770 20100 7774 20156
rect 7774 20100 7830 20156
rect 7830 20100 7834 20156
rect 7770 20096 7834 20100
rect 7850 20156 7914 20160
rect 7850 20100 7854 20156
rect 7854 20100 7910 20156
rect 7910 20100 7914 20156
rect 7850 20096 7914 20100
rect 12049 20156 12113 20160
rect 12049 20100 12053 20156
rect 12053 20100 12109 20156
rect 12109 20100 12113 20156
rect 12049 20096 12113 20100
rect 12129 20156 12193 20160
rect 12129 20100 12133 20156
rect 12133 20100 12189 20156
rect 12189 20100 12193 20156
rect 12129 20096 12193 20100
rect 12209 20156 12273 20160
rect 12209 20100 12213 20156
rect 12213 20100 12269 20156
rect 12269 20100 12273 20156
rect 12209 20096 12273 20100
rect 12289 20156 12353 20160
rect 12289 20100 12293 20156
rect 12293 20100 12349 20156
rect 12349 20100 12353 20156
rect 12289 20096 12353 20100
rect 16488 20156 16552 20160
rect 16488 20100 16492 20156
rect 16492 20100 16548 20156
rect 16548 20100 16552 20156
rect 16488 20096 16552 20100
rect 16568 20156 16632 20160
rect 16568 20100 16572 20156
rect 16572 20100 16628 20156
rect 16628 20100 16632 20156
rect 16568 20096 16632 20100
rect 16648 20156 16712 20160
rect 16648 20100 16652 20156
rect 16652 20100 16708 20156
rect 16708 20100 16712 20156
rect 16648 20096 16712 20100
rect 16728 20156 16792 20160
rect 16728 20100 16732 20156
rect 16732 20100 16788 20156
rect 16788 20100 16792 20156
rect 16728 20096 16792 20100
rect 5390 19612 5454 19616
rect 5390 19556 5394 19612
rect 5394 19556 5450 19612
rect 5450 19556 5454 19612
rect 5390 19552 5454 19556
rect 5470 19612 5534 19616
rect 5470 19556 5474 19612
rect 5474 19556 5530 19612
rect 5530 19556 5534 19612
rect 5470 19552 5534 19556
rect 5550 19612 5614 19616
rect 5550 19556 5554 19612
rect 5554 19556 5610 19612
rect 5610 19556 5614 19612
rect 5550 19552 5614 19556
rect 5630 19612 5694 19616
rect 5630 19556 5634 19612
rect 5634 19556 5690 19612
rect 5690 19556 5694 19612
rect 5630 19552 5694 19556
rect 9829 19612 9893 19616
rect 9829 19556 9833 19612
rect 9833 19556 9889 19612
rect 9889 19556 9893 19612
rect 9829 19552 9893 19556
rect 9909 19612 9973 19616
rect 9909 19556 9913 19612
rect 9913 19556 9969 19612
rect 9969 19556 9973 19612
rect 9909 19552 9973 19556
rect 9989 19612 10053 19616
rect 9989 19556 9993 19612
rect 9993 19556 10049 19612
rect 10049 19556 10053 19612
rect 9989 19552 10053 19556
rect 10069 19612 10133 19616
rect 10069 19556 10073 19612
rect 10073 19556 10129 19612
rect 10129 19556 10133 19612
rect 10069 19552 10133 19556
rect 14268 19612 14332 19616
rect 14268 19556 14272 19612
rect 14272 19556 14328 19612
rect 14328 19556 14332 19612
rect 14268 19552 14332 19556
rect 14348 19612 14412 19616
rect 14348 19556 14352 19612
rect 14352 19556 14408 19612
rect 14408 19556 14412 19612
rect 14348 19552 14412 19556
rect 14428 19612 14492 19616
rect 14428 19556 14432 19612
rect 14432 19556 14488 19612
rect 14488 19556 14492 19612
rect 14428 19552 14492 19556
rect 14508 19612 14572 19616
rect 14508 19556 14512 19612
rect 14512 19556 14568 19612
rect 14568 19556 14572 19612
rect 14508 19552 14572 19556
rect 18707 19612 18771 19616
rect 18707 19556 18711 19612
rect 18711 19556 18767 19612
rect 18767 19556 18771 19612
rect 18707 19552 18771 19556
rect 18787 19612 18851 19616
rect 18787 19556 18791 19612
rect 18791 19556 18847 19612
rect 18847 19556 18851 19612
rect 18787 19552 18851 19556
rect 18867 19612 18931 19616
rect 18867 19556 18871 19612
rect 18871 19556 18927 19612
rect 18927 19556 18931 19612
rect 18867 19552 18931 19556
rect 18947 19612 19011 19616
rect 18947 19556 18951 19612
rect 18951 19556 19007 19612
rect 19007 19556 19011 19612
rect 18947 19552 19011 19556
rect 3171 19068 3235 19072
rect 3171 19012 3175 19068
rect 3175 19012 3231 19068
rect 3231 19012 3235 19068
rect 3171 19008 3235 19012
rect 3251 19068 3315 19072
rect 3251 19012 3255 19068
rect 3255 19012 3311 19068
rect 3311 19012 3315 19068
rect 3251 19008 3315 19012
rect 3331 19068 3395 19072
rect 3331 19012 3335 19068
rect 3335 19012 3391 19068
rect 3391 19012 3395 19068
rect 3331 19008 3395 19012
rect 3411 19068 3475 19072
rect 3411 19012 3415 19068
rect 3415 19012 3471 19068
rect 3471 19012 3475 19068
rect 3411 19008 3475 19012
rect 7610 19068 7674 19072
rect 7610 19012 7614 19068
rect 7614 19012 7670 19068
rect 7670 19012 7674 19068
rect 7610 19008 7674 19012
rect 7690 19068 7754 19072
rect 7690 19012 7694 19068
rect 7694 19012 7750 19068
rect 7750 19012 7754 19068
rect 7690 19008 7754 19012
rect 7770 19068 7834 19072
rect 7770 19012 7774 19068
rect 7774 19012 7830 19068
rect 7830 19012 7834 19068
rect 7770 19008 7834 19012
rect 7850 19068 7914 19072
rect 7850 19012 7854 19068
rect 7854 19012 7910 19068
rect 7910 19012 7914 19068
rect 7850 19008 7914 19012
rect 12049 19068 12113 19072
rect 12049 19012 12053 19068
rect 12053 19012 12109 19068
rect 12109 19012 12113 19068
rect 12049 19008 12113 19012
rect 12129 19068 12193 19072
rect 12129 19012 12133 19068
rect 12133 19012 12189 19068
rect 12189 19012 12193 19068
rect 12129 19008 12193 19012
rect 12209 19068 12273 19072
rect 12209 19012 12213 19068
rect 12213 19012 12269 19068
rect 12269 19012 12273 19068
rect 12209 19008 12273 19012
rect 12289 19068 12353 19072
rect 12289 19012 12293 19068
rect 12293 19012 12349 19068
rect 12349 19012 12353 19068
rect 12289 19008 12353 19012
rect 16488 19068 16552 19072
rect 16488 19012 16492 19068
rect 16492 19012 16548 19068
rect 16548 19012 16552 19068
rect 16488 19008 16552 19012
rect 16568 19068 16632 19072
rect 16568 19012 16572 19068
rect 16572 19012 16628 19068
rect 16628 19012 16632 19068
rect 16568 19008 16632 19012
rect 16648 19068 16712 19072
rect 16648 19012 16652 19068
rect 16652 19012 16708 19068
rect 16708 19012 16712 19068
rect 16648 19008 16712 19012
rect 16728 19068 16792 19072
rect 16728 19012 16732 19068
rect 16732 19012 16788 19068
rect 16788 19012 16792 19068
rect 16728 19008 16792 19012
rect 5390 18524 5454 18528
rect 5390 18468 5394 18524
rect 5394 18468 5450 18524
rect 5450 18468 5454 18524
rect 5390 18464 5454 18468
rect 5470 18524 5534 18528
rect 5470 18468 5474 18524
rect 5474 18468 5530 18524
rect 5530 18468 5534 18524
rect 5470 18464 5534 18468
rect 5550 18524 5614 18528
rect 5550 18468 5554 18524
rect 5554 18468 5610 18524
rect 5610 18468 5614 18524
rect 5550 18464 5614 18468
rect 5630 18524 5694 18528
rect 5630 18468 5634 18524
rect 5634 18468 5690 18524
rect 5690 18468 5694 18524
rect 5630 18464 5694 18468
rect 9829 18524 9893 18528
rect 9829 18468 9833 18524
rect 9833 18468 9889 18524
rect 9889 18468 9893 18524
rect 9829 18464 9893 18468
rect 9909 18524 9973 18528
rect 9909 18468 9913 18524
rect 9913 18468 9969 18524
rect 9969 18468 9973 18524
rect 9909 18464 9973 18468
rect 9989 18524 10053 18528
rect 9989 18468 9993 18524
rect 9993 18468 10049 18524
rect 10049 18468 10053 18524
rect 9989 18464 10053 18468
rect 10069 18524 10133 18528
rect 10069 18468 10073 18524
rect 10073 18468 10129 18524
rect 10129 18468 10133 18524
rect 10069 18464 10133 18468
rect 14268 18524 14332 18528
rect 14268 18468 14272 18524
rect 14272 18468 14328 18524
rect 14328 18468 14332 18524
rect 14268 18464 14332 18468
rect 14348 18524 14412 18528
rect 14348 18468 14352 18524
rect 14352 18468 14408 18524
rect 14408 18468 14412 18524
rect 14348 18464 14412 18468
rect 14428 18524 14492 18528
rect 14428 18468 14432 18524
rect 14432 18468 14488 18524
rect 14488 18468 14492 18524
rect 14428 18464 14492 18468
rect 14508 18524 14572 18528
rect 14508 18468 14512 18524
rect 14512 18468 14568 18524
rect 14568 18468 14572 18524
rect 14508 18464 14572 18468
rect 18707 18524 18771 18528
rect 18707 18468 18711 18524
rect 18711 18468 18767 18524
rect 18767 18468 18771 18524
rect 18707 18464 18771 18468
rect 18787 18524 18851 18528
rect 18787 18468 18791 18524
rect 18791 18468 18847 18524
rect 18847 18468 18851 18524
rect 18787 18464 18851 18468
rect 18867 18524 18931 18528
rect 18867 18468 18871 18524
rect 18871 18468 18927 18524
rect 18927 18468 18931 18524
rect 18867 18464 18931 18468
rect 18947 18524 19011 18528
rect 18947 18468 18951 18524
rect 18951 18468 19007 18524
rect 19007 18468 19011 18524
rect 18947 18464 19011 18468
rect 3171 17980 3235 17984
rect 3171 17924 3175 17980
rect 3175 17924 3231 17980
rect 3231 17924 3235 17980
rect 3171 17920 3235 17924
rect 3251 17980 3315 17984
rect 3251 17924 3255 17980
rect 3255 17924 3311 17980
rect 3311 17924 3315 17980
rect 3251 17920 3315 17924
rect 3331 17980 3395 17984
rect 3331 17924 3335 17980
rect 3335 17924 3391 17980
rect 3391 17924 3395 17980
rect 3331 17920 3395 17924
rect 3411 17980 3475 17984
rect 3411 17924 3415 17980
rect 3415 17924 3471 17980
rect 3471 17924 3475 17980
rect 3411 17920 3475 17924
rect 7610 17980 7674 17984
rect 7610 17924 7614 17980
rect 7614 17924 7670 17980
rect 7670 17924 7674 17980
rect 7610 17920 7674 17924
rect 7690 17980 7754 17984
rect 7690 17924 7694 17980
rect 7694 17924 7750 17980
rect 7750 17924 7754 17980
rect 7690 17920 7754 17924
rect 7770 17980 7834 17984
rect 7770 17924 7774 17980
rect 7774 17924 7830 17980
rect 7830 17924 7834 17980
rect 7770 17920 7834 17924
rect 7850 17980 7914 17984
rect 7850 17924 7854 17980
rect 7854 17924 7910 17980
rect 7910 17924 7914 17980
rect 7850 17920 7914 17924
rect 12049 17980 12113 17984
rect 12049 17924 12053 17980
rect 12053 17924 12109 17980
rect 12109 17924 12113 17980
rect 12049 17920 12113 17924
rect 12129 17980 12193 17984
rect 12129 17924 12133 17980
rect 12133 17924 12189 17980
rect 12189 17924 12193 17980
rect 12129 17920 12193 17924
rect 12209 17980 12273 17984
rect 12209 17924 12213 17980
rect 12213 17924 12269 17980
rect 12269 17924 12273 17980
rect 12209 17920 12273 17924
rect 12289 17980 12353 17984
rect 12289 17924 12293 17980
rect 12293 17924 12349 17980
rect 12349 17924 12353 17980
rect 12289 17920 12353 17924
rect 16488 17980 16552 17984
rect 16488 17924 16492 17980
rect 16492 17924 16548 17980
rect 16548 17924 16552 17980
rect 16488 17920 16552 17924
rect 16568 17980 16632 17984
rect 16568 17924 16572 17980
rect 16572 17924 16628 17980
rect 16628 17924 16632 17980
rect 16568 17920 16632 17924
rect 16648 17980 16712 17984
rect 16648 17924 16652 17980
rect 16652 17924 16708 17980
rect 16708 17924 16712 17980
rect 16648 17920 16712 17924
rect 16728 17980 16792 17984
rect 16728 17924 16732 17980
rect 16732 17924 16788 17980
rect 16788 17924 16792 17980
rect 16728 17920 16792 17924
rect 5390 17436 5454 17440
rect 5390 17380 5394 17436
rect 5394 17380 5450 17436
rect 5450 17380 5454 17436
rect 5390 17376 5454 17380
rect 5470 17436 5534 17440
rect 5470 17380 5474 17436
rect 5474 17380 5530 17436
rect 5530 17380 5534 17436
rect 5470 17376 5534 17380
rect 5550 17436 5614 17440
rect 5550 17380 5554 17436
rect 5554 17380 5610 17436
rect 5610 17380 5614 17436
rect 5550 17376 5614 17380
rect 5630 17436 5694 17440
rect 5630 17380 5634 17436
rect 5634 17380 5690 17436
rect 5690 17380 5694 17436
rect 5630 17376 5694 17380
rect 9829 17436 9893 17440
rect 9829 17380 9833 17436
rect 9833 17380 9889 17436
rect 9889 17380 9893 17436
rect 9829 17376 9893 17380
rect 9909 17436 9973 17440
rect 9909 17380 9913 17436
rect 9913 17380 9969 17436
rect 9969 17380 9973 17436
rect 9909 17376 9973 17380
rect 9989 17436 10053 17440
rect 9989 17380 9993 17436
rect 9993 17380 10049 17436
rect 10049 17380 10053 17436
rect 9989 17376 10053 17380
rect 10069 17436 10133 17440
rect 10069 17380 10073 17436
rect 10073 17380 10129 17436
rect 10129 17380 10133 17436
rect 10069 17376 10133 17380
rect 14268 17436 14332 17440
rect 14268 17380 14272 17436
rect 14272 17380 14328 17436
rect 14328 17380 14332 17436
rect 14268 17376 14332 17380
rect 14348 17436 14412 17440
rect 14348 17380 14352 17436
rect 14352 17380 14408 17436
rect 14408 17380 14412 17436
rect 14348 17376 14412 17380
rect 14428 17436 14492 17440
rect 14428 17380 14432 17436
rect 14432 17380 14488 17436
rect 14488 17380 14492 17436
rect 14428 17376 14492 17380
rect 14508 17436 14572 17440
rect 14508 17380 14512 17436
rect 14512 17380 14568 17436
rect 14568 17380 14572 17436
rect 14508 17376 14572 17380
rect 18707 17436 18771 17440
rect 18707 17380 18711 17436
rect 18711 17380 18767 17436
rect 18767 17380 18771 17436
rect 18707 17376 18771 17380
rect 18787 17436 18851 17440
rect 18787 17380 18791 17436
rect 18791 17380 18847 17436
rect 18847 17380 18851 17436
rect 18787 17376 18851 17380
rect 18867 17436 18931 17440
rect 18867 17380 18871 17436
rect 18871 17380 18927 17436
rect 18927 17380 18931 17436
rect 18867 17376 18931 17380
rect 18947 17436 19011 17440
rect 18947 17380 18951 17436
rect 18951 17380 19007 17436
rect 19007 17380 19011 17436
rect 18947 17376 19011 17380
rect 3171 16892 3235 16896
rect 3171 16836 3175 16892
rect 3175 16836 3231 16892
rect 3231 16836 3235 16892
rect 3171 16832 3235 16836
rect 3251 16892 3315 16896
rect 3251 16836 3255 16892
rect 3255 16836 3311 16892
rect 3311 16836 3315 16892
rect 3251 16832 3315 16836
rect 3331 16892 3395 16896
rect 3331 16836 3335 16892
rect 3335 16836 3391 16892
rect 3391 16836 3395 16892
rect 3331 16832 3395 16836
rect 3411 16892 3475 16896
rect 3411 16836 3415 16892
rect 3415 16836 3471 16892
rect 3471 16836 3475 16892
rect 3411 16832 3475 16836
rect 7610 16892 7674 16896
rect 7610 16836 7614 16892
rect 7614 16836 7670 16892
rect 7670 16836 7674 16892
rect 7610 16832 7674 16836
rect 7690 16892 7754 16896
rect 7690 16836 7694 16892
rect 7694 16836 7750 16892
rect 7750 16836 7754 16892
rect 7690 16832 7754 16836
rect 7770 16892 7834 16896
rect 7770 16836 7774 16892
rect 7774 16836 7830 16892
rect 7830 16836 7834 16892
rect 7770 16832 7834 16836
rect 7850 16892 7914 16896
rect 7850 16836 7854 16892
rect 7854 16836 7910 16892
rect 7910 16836 7914 16892
rect 7850 16832 7914 16836
rect 12049 16892 12113 16896
rect 12049 16836 12053 16892
rect 12053 16836 12109 16892
rect 12109 16836 12113 16892
rect 12049 16832 12113 16836
rect 12129 16892 12193 16896
rect 12129 16836 12133 16892
rect 12133 16836 12189 16892
rect 12189 16836 12193 16892
rect 12129 16832 12193 16836
rect 12209 16892 12273 16896
rect 12209 16836 12213 16892
rect 12213 16836 12269 16892
rect 12269 16836 12273 16892
rect 12209 16832 12273 16836
rect 12289 16892 12353 16896
rect 12289 16836 12293 16892
rect 12293 16836 12349 16892
rect 12349 16836 12353 16892
rect 12289 16832 12353 16836
rect 16488 16892 16552 16896
rect 16488 16836 16492 16892
rect 16492 16836 16548 16892
rect 16548 16836 16552 16892
rect 16488 16832 16552 16836
rect 16568 16892 16632 16896
rect 16568 16836 16572 16892
rect 16572 16836 16628 16892
rect 16628 16836 16632 16892
rect 16568 16832 16632 16836
rect 16648 16892 16712 16896
rect 16648 16836 16652 16892
rect 16652 16836 16708 16892
rect 16708 16836 16712 16892
rect 16648 16832 16712 16836
rect 16728 16892 16792 16896
rect 16728 16836 16732 16892
rect 16732 16836 16788 16892
rect 16788 16836 16792 16892
rect 16728 16832 16792 16836
rect 5390 16348 5454 16352
rect 5390 16292 5394 16348
rect 5394 16292 5450 16348
rect 5450 16292 5454 16348
rect 5390 16288 5454 16292
rect 5470 16348 5534 16352
rect 5470 16292 5474 16348
rect 5474 16292 5530 16348
rect 5530 16292 5534 16348
rect 5470 16288 5534 16292
rect 5550 16348 5614 16352
rect 5550 16292 5554 16348
rect 5554 16292 5610 16348
rect 5610 16292 5614 16348
rect 5550 16288 5614 16292
rect 5630 16348 5694 16352
rect 5630 16292 5634 16348
rect 5634 16292 5690 16348
rect 5690 16292 5694 16348
rect 5630 16288 5694 16292
rect 9829 16348 9893 16352
rect 9829 16292 9833 16348
rect 9833 16292 9889 16348
rect 9889 16292 9893 16348
rect 9829 16288 9893 16292
rect 9909 16348 9973 16352
rect 9909 16292 9913 16348
rect 9913 16292 9969 16348
rect 9969 16292 9973 16348
rect 9909 16288 9973 16292
rect 9989 16348 10053 16352
rect 9989 16292 9993 16348
rect 9993 16292 10049 16348
rect 10049 16292 10053 16348
rect 9989 16288 10053 16292
rect 10069 16348 10133 16352
rect 10069 16292 10073 16348
rect 10073 16292 10129 16348
rect 10129 16292 10133 16348
rect 10069 16288 10133 16292
rect 14268 16348 14332 16352
rect 14268 16292 14272 16348
rect 14272 16292 14328 16348
rect 14328 16292 14332 16348
rect 14268 16288 14332 16292
rect 14348 16348 14412 16352
rect 14348 16292 14352 16348
rect 14352 16292 14408 16348
rect 14408 16292 14412 16348
rect 14348 16288 14412 16292
rect 14428 16348 14492 16352
rect 14428 16292 14432 16348
rect 14432 16292 14488 16348
rect 14488 16292 14492 16348
rect 14428 16288 14492 16292
rect 14508 16348 14572 16352
rect 14508 16292 14512 16348
rect 14512 16292 14568 16348
rect 14568 16292 14572 16348
rect 14508 16288 14572 16292
rect 18707 16348 18771 16352
rect 18707 16292 18711 16348
rect 18711 16292 18767 16348
rect 18767 16292 18771 16348
rect 18707 16288 18771 16292
rect 18787 16348 18851 16352
rect 18787 16292 18791 16348
rect 18791 16292 18847 16348
rect 18847 16292 18851 16348
rect 18787 16288 18851 16292
rect 18867 16348 18931 16352
rect 18867 16292 18871 16348
rect 18871 16292 18927 16348
rect 18927 16292 18931 16348
rect 18867 16288 18931 16292
rect 18947 16348 19011 16352
rect 18947 16292 18951 16348
rect 18951 16292 19007 16348
rect 19007 16292 19011 16348
rect 18947 16288 19011 16292
rect 3171 15804 3235 15808
rect 3171 15748 3175 15804
rect 3175 15748 3231 15804
rect 3231 15748 3235 15804
rect 3171 15744 3235 15748
rect 3251 15804 3315 15808
rect 3251 15748 3255 15804
rect 3255 15748 3311 15804
rect 3311 15748 3315 15804
rect 3251 15744 3315 15748
rect 3331 15804 3395 15808
rect 3331 15748 3335 15804
rect 3335 15748 3391 15804
rect 3391 15748 3395 15804
rect 3331 15744 3395 15748
rect 3411 15804 3475 15808
rect 3411 15748 3415 15804
rect 3415 15748 3471 15804
rect 3471 15748 3475 15804
rect 3411 15744 3475 15748
rect 7610 15804 7674 15808
rect 7610 15748 7614 15804
rect 7614 15748 7670 15804
rect 7670 15748 7674 15804
rect 7610 15744 7674 15748
rect 7690 15804 7754 15808
rect 7690 15748 7694 15804
rect 7694 15748 7750 15804
rect 7750 15748 7754 15804
rect 7690 15744 7754 15748
rect 7770 15804 7834 15808
rect 7770 15748 7774 15804
rect 7774 15748 7830 15804
rect 7830 15748 7834 15804
rect 7770 15744 7834 15748
rect 7850 15804 7914 15808
rect 7850 15748 7854 15804
rect 7854 15748 7910 15804
rect 7910 15748 7914 15804
rect 7850 15744 7914 15748
rect 12049 15804 12113 15808
rect 12049 15748 12053 15804
rect 12053 15748 12109 15804
rect 12109 15748 12113 15804
rect 12049 15744 12113 15748
rect 12129 15804 12193 15808
rect 12129 15748 12133 15804
rect 12133 15748 12189 15804
rect 12189 15748 12193 15804
rect 12129 15744 12193 15748
rect 12209 15804 12273 15808
rect 12209 15748 12213 15804
rect 12213 15748 12269 15804
rect 12269 15748 12273 15804
rect 12209 15744 12273 15748
rect 12289 15804 12353 15808
rect 12289 15748 12293 15804
rect 12293 15748 12349 15804
rect 12349 15748 12353 15804
rect 12289 15744 12353 15748
rect 16488 15804 16552 15808
rect 16488 15748 16492 15804
rect 16492 15748 16548 15804
rect 16548 15748 16552 15804
rect 16488 15744 16552 15748
rect 16568 15804 16632 15808
rect 16568 15748 16572 15804
rect 16572 15748 16628 15804
rect 16628 15748 16632 15804
rect 16568 15744 16632 15748
rect 16648 15804 16712 15808
rect 16648 15748 16652 15804
rect 16652 15748 16708 15804
rect 16708 15748 16712 15804
rect 16648 15744 16712 15748
rect 16728 15804 16792 15808
rect 16728 15748 16732 15804
rect 16732 15748 16788 15804
rect 16788 15748 16792 15804
rect 16728 15744 16792 15748
rect 5390 15260 5454 15264
rect 5390 15204 5394 15260
rect 5394 15204 5450 15260
rect 5450 15204 5454 15260
rect 5390 15200 5454 15204
rect 5470 15260 5534 15264
rect 5470 15204 5474 15260
rect 5474 15204 5530 15260
rect 5530 15204 5534 15260
rect 5470 15200 5534 15204
rect 5550 15260 5614 15264
rect 5550 15204 5554 15260
rect 5554 15204 5610 15260
rect 5610 15204 5614 15260
rect 5550 15200 5614 15204
rect 5630 15260 5694 15264
rect 5630 15204 5634 15260
rect 5634 15204 5690 15260
rect 5690 15204 5694 15260
rect 5630 15200 5694 15204
rect 9829 15260 9893 15264
rect 9829 15204 9833 15260
rect 9833 15204 9889 15260
rect 9889 15204 9893 15260
rect 9829 15200 9893 15204
rect 9909 15260 9973 15264
rect 9909 15204 9913 15260
rect 9913 15204 9969 15260
rect 9969 15204 9973 15260
rect 9909 15200 9973 15204
rect 9989 15260 10053 15264
rect 9989 15204 9993 15260
rect 9993 15204 10049 15260
rect 10049 15204 10053 15260
rect 9989 15200 10053 15204
rect 10069 15260 10133 15264
rect 10069 15204 10073 15260
rect 10073 15204 10129 15260
rect 10129 15204 10133 15260
rect 10069 15200 10133 15204
rect 14268 15260 14332 15264
rect 14268 15204 14272 15260
rect 14272 15204 14328 15260
rect 14328 15204 14332 15260
rect 14268 15200 14332 15204
rect 14348 15260 14412 15264
rect 14348 15204 14352 15260
rect 14352 15204 14408 15260
rect 14408 15204 14412 15260
rect 14348 15200 14412 15204
rect 14428 15260 14492 15264
rect 14428 15204 14432 15260
rect 14432 15204 14488 15260
rect 14488 15204 14492 15260
rect 14428 15200 14492 15204
rect 14508 15260 14572 15264
rect 14508 15204 14512 15260
rect 14512 15204 14568 15260
rect 14568 15204 14572 15260
rect 14508 15200 14572 15204
rect 18707 15260 18771 15264
rect 18707 15204 18711 15260
rect 18711 15204 18767 15260
rect 18767 15204 18771 15260
rect 18707 15200 18771 15204
rect 18787 15260 18851 15264
rect 18787 15204 18791 15260
rect 18791 15204 18847 15260
rect 18847 15204 18851 15260
rect 18787 15200 18851 15204
rect 18867 15260 18931 15264
rect 18867 15204 18871 15260
rect 18871 15204 18927 15260
rect 18927 15204 18931 15260
rect 18867 15200 18931 15204
rect 18947 15260 19011 15264
rect 18947 15204 18951 15260
rect 18951 15204 19007 15260
rect 19007 15204 19011 15260
rect 18947 15200 19011 15204
rect 3171 14716 3235 14720
rect 3171 14660 3175 14716
rect 3175 14660 3231 14716
rect 3231 14660 3235 14716
rect 3171 14656 3235 14660
rect 3251 14716 3315 14720
rect 3251 14660 3255 14716
rect 3255 14660 3311 14716
rect 3311 14660 3315 14716
rect 3251 14656 3315 14660
rect 3331 14716 3395 14720
rect 3331 14660 3335 14716
rect 3335 14660 3391 14716
rect 3391 14660 3395 14716
rect 3331 14656 3395 14660
rect 3411 14716 3475 14720
rect 3411 14660 3415 14716
rect 3415 14660 3471 14716
rect 3471 14660 3475 14716
rect 3411 14656 3475 14660
rect 7610 14716 7674 14720
rect 7610 14660 7614 14716
rect 7614 14660 7670 14716
rect 7670 14660 7674 14716
rect 7610 14656 7674 14660
rect 7690 14716 7754 14720
rect 7690 14660 7694 14716
rect 7694 14660 7750 14716
rect 7750 14660 7754 14716
rect 7690 14656 7754 14660
rect 7770 14716 7834 14720
rect 7770 14660 7774 14716
rect 7774 14660 7830 14716
rect 7830 14660 7834 14716
rect 7770 14656 7834 14660
rect 7850 14716 7914 14720
rect 7850 14660 7854 14716
rect 7854 14660 7910 14716
rect 7910 14660 7914 14716
rect 7850 14656 7914 14660
rect 12049 14716 12113 14720
rect 12049 14660 12053 14716
rect 12053 14660 12109 14716
rect 12109 14660 12113 14716
rect 12049 14656 12113 14660
rect 12129 14716 12193 14720
rect 12129 14660 12133 14716
rect 12133 14660 12189 14716
rect 12189 14660 12193 14716
rect 12129 14656 12193 14660
rect 12209 14716 12273 14720
rect 12209 14660 12213 14716
rect 12213 14660 12269 14716
rect 12269 14660 12273 14716
rect 12209 14656 12273 14660
rect 12289 14716 12353 14720
rect 12289 14660 12293 14716
rect 12293 14660 12349 14716
rect 12349 14660 12353 14716
rect 12289 14656 12353 14660
rect 16488 14716 16552 14720
rect 16488 14660 16492 14716
rect 16492 14660 16548 14716
rect 16548 14660 16552 14716
rect 16488 14656 16552 14660
rect 16568 14716 16632 14720
rect 16568 14660 16572 14716
rect 16572 14660 16628 14716
rect 16628 14660 16632 14716
rect 16568 14656 16632 14660
rect 16648 14716 16712 14720
rect 16648 14660 16652 14716
rect 16652 14660 16708 14716
rect 16708 14660 16712 14716
rect 16648 14656 16712 14660
rect 16728 14716 16792 14720
rect 16728 14660 16732 14716
rect 16732 14660 16788 14716
rect 16788 14660 16792 14716
rect 16728 14656 16792 14660
rect 5390 14172 5454 14176
rect 5390 14116 5394 14172
rect 5394 14116 5450 14172
rect 5450 14116 5454 14172
rect 5390 14112 5454 14116
rect 5470 14172 5534 14176
rect 5470 14116 5474 14172
rect 5474 14116 5530 14172
rect 5530 14116 5534 14172
rect 5470 14112 5534 14116
rect 5550 14172 5614 14176
rect 5550 14116 5554 14172
rect 5554 14116 5610 14172
rect 5610 14116 5614 14172
rect 5550 14112 5614 14116
rect 5630 14172 5694 14176
rect 5630 14116 5634 14172
rect 5634 14116 5690 14172
rect 5690 14116 5694 14172
rect 5630 14112 5694 14116
rect 9829 14172 9893 14176
rect 9829 14116 9833 14172
rect 9833 14116 9889 14172
rect 9889 14116 9893 14172
rect 9829 14112 9893 14116
rect 9909 14172 9973 14176
rect 9909 14116 9913 14172
rect 9913 14116 9969 14172
rect 9969 14116 9973 14172
rect 9909 14112 9973 14116
rect 9989 14172 10053 14176
rect 9989 14116 9993 14172
rect 9993 14116 10049 14172
rect 10049 14116 10053 14172
rect 9989 14112 10053 14116
rect 10069 14172 10133 14176
rect 10069 14116 10073 14172
rect 10073 14116 10129 14172
rect 10129 14116 10133 14172
rect 10069 14112 10133 14116
rect 14268 14172 14332 14176
rect 14268 14116 14272 14172
rect 14272 14116 14328 14172
rect 14328 14116 14332 14172
rect 14268 14112 14332 14116
rect 14348 14172 14412 14176
rect 14348 14116 14352 14172
rect 14352 14116 14408 14172
rect 14408 14116 14412 14172
rect 14348 14112 14412 14116
rect 14428 14172 14492 14176
rect 14428 14116 14432 14172
rect 14432 14116 14488 14172
rect 14488 14116 14492 14172
rect 14428 14112 14492 14116
rect 14508 14172 14572 14176
rect 14508 14116 14512 14172
rect 14512 14116 14568 14172
rect 14568 14116 14572 14172
rect 14508 14112 14572 14116
rect 18707 14172 18771 14176
rect 18707 14116 18711 14172
rect 18711 14116 18767 14172
rect 18767 14116 18771 14172
rect 18707 14112 18771 14116
rect 18787 14172 18851 14176
rect 18787 14116 18791 14172
rect 18791 14116 18847 14172
rect 18847 14116 18851 14172
rect 18787 14112 18851 14116
rect 18867 14172 18931 14176
rect 18867 14116 18871 14172
rect 18871 14116 18927 14172
rect 18927 14116 18931 14172
rect 18867 14112 18931 14116
rect 18947 14172 19011 14176
rect 18947 14116 18951 14172
rect 18951 14116 19007 14172
rect 19007 14116 19011 14172
rect 18947 14112 19011 14116
rect 3171 13628 3235 13632
rect 3171 13572 3175 13628
rect 3175 13572 3231 13628
rect 3231 13572 3235 13628
rect 3171 13568 3235 13572
rect 3251 13628 3315 13632
rect 3251 13572 3255 13628
rect 3255 13572 3311 13628
rect 3311 13572 3315 13628
rect 3251 13568 3315 13572
rect 3331 13628 3395 13632
rect 3331 13572 3335 13628
rect 3335 13572 3391 13628
rect 3391 13572 3395 13628
rect 3331 13568 3395 13572
rect 3411 13628 3475 13632
rect 3411 13572 3415 13628
rect 3415 13572 3471 13628
rect 3471 13572 3475 13628
rect 3411 13568 3475 13572
rect 7610 13628 7674 13632
rect 7610 13572 7614 13628
rect 7614 13572 7670 13628
rect 7670 13572 7674 13628
rect 7610 13568 7674 13572
rect 7690 13628 7754 13632
rect 7690 13572 7694 13628
rect 7694 13572 7750 13628
rect 7750 13572 7754 13628
rect 7690 13568 7754 13572
rect 7770 13628 7834 13632
rect 7770 13572 7774 13628
rect 7774 13572 7830 13628
rect 7830 13572 7834 13628
rect 7770 13568 7834 13572
rect 7850 13628 7914 13632
rect 7850 13572 7854 13628
rect 7854 13572 7910 13628
rect 7910 13572 7914 13628
rect 7850 13568 7914 13572
rect 12049 13628 12113 13632
rect 12049 13572 12053 13628
rect 12053 13572 12109 13628
rect 12109 13572 12113 13628
rect 12049 13568 12113 13572
rect 12129 13628 12193 13632
rect 12129 13572 12133 13628
rect 12133 13572 12189 13628
rect 12189 13572 12193 13628
rect 12129 13568 12193 13572
rect 12209 13628 12273 13632
rect 12209 13572 12213 13628
rect 12213 13572 12269 13628
rect 12269 13572 12273 13628
rect 12209 13568 12273 13572
rect 12289 13628 12353 13632
rect 12289 13572 12293 13628
rect 12293 13572 12349 13628
rect 12349 13572 12353 13628
rect 12289 13568 12353 13572
rect 16488 13628 16552 13632
rect 16488 13572 16492 13628
rect 16492 13572 16548 13628
rect 16548 13572 16552 13628
rect 16488 13568 16552 13572
rect 16568 13628 16632 13632
rect 16568 13572 16572 13628
rect 16572 13572 16628 13628
rect 16628 13572 16632 13628
rect 16568 13568 16632 13572
rect 16648 13628 16712 13632
rect 16648 13572 16652 13628
rect 16652 13572 16708 13628
rect 16708 13572 16712 13628
rect 16648 13568 16712 13572
rect 16728 13628 16792 13632
rect 16728 13572 16732 13628
rect 16732 13572 16788 13628
rect 16788 13572 16792 13628
rect 16728 13568 16792 13572
rect 5390 13084 5454 13088
rect 5390 13028 5394 13084
rect 5394 13028 5450 13084
rect 5450 13028 5454 13084
rect 5390 13024 5454 13028
rect 5470 13084 5534 13088
rect 5470 13028 5474 13084
rect 5474 13028 5530 13084
rect 5530 13028 5534 13084
rect 5470 13024 5534 13028
rect 5550 13084 5614 13088
rect 5550 13028 5554 13084
rect 5554 13028 5610 13084
rect 5610 13028 5614 13084
rect 5550 13024 5614 13028
rect 5630 13084 5694 13088
rect 5630 13028 5634 13084
rect 5634 13028 5690 13084
rect 5690 13028 5694 13084
rect 5630 13024 5694 13028
rect 9829 13084 9893 13088
rect 9829 13028 9833 13084
rect 9833 13028 9889 13084
rect 9889 13028 9893 13084
rect 9829 13024 9893 13028
rect 9909 13084 9973 13088
rect 9909 13028 9913 13084
rect 9913 13028 9969 13084
rect 9969 13028 9973 13084
rect 9909 13024 9973 13028
rect 9989 13084 10053 13088
rect 9989 13028 9993 13084
rect 9993 13028 10049 13084
rect 10049 13028 10053 13084
rect 9989 13024 10053 13028
rect 10069 13084 10133 13088
rect 10069 13028 10073 13084
rect 10073 13028 10129 13084
rect 10129 13028 10133 13084
rect 10069 13024 10133 13028
rect 14268 13084 14332 13088
rect 14268 13028 14272 13084
rect 14272 13028 14328 13084
rect 14328 13028 14332 13084
rect 14268 13024 14332 13028
rect 14348 13084 14412 13088
rect 14348 13028 14352 13084
rect 14352 13028 14408 13084
rect 14408 13028 14412 13084
rect 14348 13024 14412 13028
rect 14428 13084 14492 13088
rect 14428 13028 14432 13084
rect 14432 13028 14488 13084
rect 14488 13028 14492 13084
rect 14428 13024 14492 13028
rect 14508 13084 14572 13088
rect 14508 13028 14512 13084
rect 14512 13028 14568 13084
rect 14568 13028 14572 13084
rect 14508 13024 14572 13028
rect 18707 13084 18771 13088
rect 18707 13028 18711 13084
rect 18711 13028 18767 13084
rect 18767 13028 18771 13084
rect 18707 13024 18771 13028
rect 18787 13084 18851 13088
rect 18787 13028 18791 13084
rect 18791 13028 18847 13084
rect 18847 13028 18851 13084
rect 18787 13024 18851 13028
rect 18867 13084 18931 13088
rect 18867 13028 18871 13084
rect 18871 13028 18927 13084
rect 18927 13028 18931 13084
rect 18867 13024 18931 13028
rect 18947 13084 19011 13088
rect 18947 13028 18951 13084
rect 18951 13028 19007 13084
rect 19007 13028 19011 13084
rect 18947 13024 19011 13028
rect 3171 12540 3235 12544
rect 3171 12484 3175 12540
rect 3175 12484 3231 12540
rect 3231 12484 3235 12540
rect 3171 12480 3235 12484
rect 3251 12540 3315 12544
rect 3251 12484 3255 12540
rect 3255 12484 3311 12540
rect 3311 12484 3315 12540
rect 3251 12480 3315 12484
rect 3331 12540 3395 12544
rect 3331 12484 3335 12540
rect 3335 12484 3391 12540
rect 3391 12484 3395 12540
rect 3331 12480 3395 12484
rect 3411 12540 3475 12544
rect 3411 12484 3415 12540
rect 3415 12484 3471 12540
rect 3471 12484 3475 12540
rect 3411 12480 3475 12484
rect 7610 12540 7674 12544
rect 7610 12484 7614 12540
rect 7614 12484 7670 12540
rect 7670 12484 7674 12540
rect 7610 12480 7674 12484
rect 7690 12540 7754 12544
rect 7690 12484 7694 12540
rect 7694 12484 7750 12540
rect 7750 12484 7754 12540
rect 7690 12480 7754 12484
rect 7770 12540 7834 12544
rect 7770 12484 7774 12540
rect 7774 12484 7830 12540
rect 7830 12484 7834 12540
rect 7770 12480 7834 12484
rect 7850 12540 7914 12544
rect 7850 12484 7854 12540
rect 7854 12484 7910 12540
rect 7910 12484 7914 12540
rect 7850 12480 7914 12484
rect 12049 12540 12113 12544
rect 12049 12484 12053 12540
rect 12053 12484 12109 12540
rect 12109 12484 12113 12540
rect 12049 12480 12113 12484
rect 12129 12540 12193 12544
rect 12129 12484 12133 12540
rect 12133 12484 12189 12540
rect 12189 12484 12193 12540
rect 12129 12480 12193 12484
rect 12209 12540 12273 12544
rect 12209 12484 12213 12540
rect 12213 12484 12269 12540
rect 12269 12484 12273 12540
rect 12209 12480 12273 12484
rect 12289 12540 12353 12544
rect 12289 12484 12293 12540
rect 12293 12484 12349 12540
rect 12349 12484 12353 12540
rect 12289 12480 12353 12484
rect 16488 12540 16552 12544
rect 16488 12484 16492 12540
rect 16492 12484 16548 12540
rect 16548 12484 16552 12540
rect 16488 12480 16552 12484
rect 16568 12540 16632 12544
rect 16568 12484 16572 12540
rect 16572 12484 16628 12540
rect 16628 12484 16632 12540
rect 16568 12480 16632 12484
rect 16648 12540 16712 12544
rect 16648 12484 16652 12540
rect 16652 12484 16708 12540
rect 16708 12484 16712 12540
rect 16648 12480 16712 12484
rect 16728 12540 16792 12544
rect 16728 12484 16732 12540
rect 16732 12484 16788 12540
rect 16788 12484 16792 12540
rect 16728 12480 16792 12484
rect 5390 11996 5454 12000
rect 5390 11940 5394 11996
rect 5394 11940 5450 11996
rect 5450 11940 5454 11996
rect 5390 11936 5454 11940
rect 5470 11996 5534 12000
rect 5470 11940 5474 11996
rect 5474 11940 5530 11996
rect 5530 11940 5534 11996
rect 5470 11936 5534 11940
rect 5550 11996 5614 12000
rect 5550 11940 5554 11996
rect 5554 11940 5610 11996
rect 5610 11940 5614 11996
rect 5550 11936 5614 11940
rect 5630 11996 5694 12000
rect 5630 11940 5634 11996
rect 5634 11940 5690 11996
rect 5690 11940 5694 11996
rect 5630 11936 5694 11940
rect 9829 11996 9893 12000
rect 9829 11940 9833 11996
rect 9833 11940 9889 11996
rect 9889 11940 9893 11996
rect 9829 11936 9893 11940
rect 9909 11996 9973 12000
rect 9909 11940 9913 11996
rect 9913 11940 9969 11996
rect 9969 11940 9973 11996
rect 9909 11936 9973 11940
rect 9989 11996 10053 12000
rect 9989 11940 9993 11996
rect 9993 11940 10049 11996
rect 10049 11940 10053 11996
rect 9989 11936 10053 11940
rect 10069 11996 10133 12000
rect 10069 11940 10073 11996
rect 10073 11940 10129 11996
rect 10129 11940 10133 11996
rect 10069 11936 10133 11940
rect 14268 11996 14332 12000
rect 14268 11940 14272 11996
rect 14272 11940 14328 11996
rect 14328 11940 14332 11996
rect 14268 11936 14332 11940
rect 14348 11996 14412 12000
rect 14348 11940 14352 11996
rect 14352 11940 14408 11996
rect 14408 11940 14412 11996
rect 14348 11936 14412 11940
rect 14428 11996 14492 12000
rect 14428 11940 14432 11996
rect 14432 11940 14488 11996
rect 14488 11940 14492 11996
rect 14428 11936 14492 11940
rect 14508 11996 14572 12000
rect 14508 11940 14512 11996
rect 14512 11940 14568 11996
rect 14568 11940 14572 11996
rect 14508 11936 14572 11940
rect 18707 11996 18771 12000
rect 18707 11940 18711 11996
rect 18711 11940 18767 11996
rect 18767 11940 18771 11996
rect 18707 11936 18771 11940
rect 18787 11996 18851 12000
rect 18787 11940 18791 11996
rect 18791 11940 18847 11996
rect 18847 11940 18851 11996
rect 18787 11936 18851 11940
rect 18867 11996 18931 12000
rect 18867 11940 18871 11996
rect 18871 11940 18927 11996
rect 18927 11940 18931 11996
rect 18867 11936 18931 11940
rect 18947 11996 19011 12000
rect 18947 11940 18951 11996
rect 18951 11940 19007 11996
rect 19007 11940 19011 11996
rect 18947 11936 19011 11940
rect 3171 11452 3235 11456
rect 3171 11396 3175 11452
rect 3175 11396 3231 11452
rect 3231 11396 3235 11452
rect 3171 11392 3235 11396
rect 3251 11452 3315 11456
rect 3251 11396 3255 11452
rect 3255 11396 3311 11452
rect 3311 11396 3315 11452
rect 3251 11392 3315 11396
rect 3331 11452 3395 11456
rect 3331 11396 3335 11452
rect 3335 11396 3391 11452
rect 3391 11396 3395 11452
rect 3331 11392 3395 11396
rect 3411 11452 3475 11456
rect 3411 11396 3415 11452
rect 3415 11396 3471 11452
rect 3471 11396 3475 11452
rect 3411 11392 3475 11396
rect 7610 11452 7674 11456
rect 7610 11396 7614 11452
rect 7614 11396 7670 11452
rect 7670 11396 7674 11452
rect 7610 11392 7674 11396
rect 7690 11452 7754 11456
rect 7690 11396 7694 11452
rect 7694 11396 7750 11452
rect 7750 11396 7754 11452
rect 7690 11392 7754 11396
rect 7770 11452 7834 11456
rect 7770 11396 7774 11452
rect 7774 11396 7830 11452
rect 7830 11396 7834 11452
rect 7770 11392 7834 11396
rect 7850 11452 7914 11456
rect 7850 11396 7854 11452
rect 7854 11396 7910 11452
rect 7910 11396 7914 11452
rect 7850 11392 7914 11396
rect 12049 11452 12113 11456
rect 12049 11396 12053 11452
rect 12053 11396 12109 11452
rect 12109 11396 12113 11452
rect 12049 11392 12113 11396
rect 12129 11452 12193 11456
rect 12129 11396 12133 11452
rect 12133 11396 12189 11452
rect 12189 11396 12193 11452
rect 12129 11392 12193 11396
rect 12209 11452 12273 11456
rect 12209 11396 12213 11452
rect 12213 11396 12269 11452
rect 12269 11396 12273 11452
rect 12209 11392 12273 11396
rect 12289 11452 12353 11456
rect 12289 11396 12293 11452
rect 12293 11396 12349 11452
rect 12349 11396 12353 11452
rect 12289 11392 12353 11396
rect 16488 11452 16552 11456
rect 16488 11396 16492 11452
rect 16492 11396 16548 11452
rect 16548 11396 16552 11452
rect 16488 11392 16552 11396
rect 16568 11452 16632 11456
rect 16568 11396 16572 11452
rect 16572 11396 16628 11452
rect 16628 11396 16632 11452
rect 16568 11392 16632 11396
rect 16648 11452 16712 11456
rect 16648 11396 16652 11452
rect 16652 11396 16708 11452
rect 16708 11396 16712 11452
rect 16648 11392 16712 11396
rect 16728 11452 16792 11456
rect 16728 11396 16732 11452
rect 16732 11396 16788 11452
rect 16788 11396 16792 11452
rect 16728 11392 16792 11396
rect 5390 10908 5454 10912
rect 5390 10852 5394 10908
rect 5394 10852 5450 10908
rect 5450 10852 5454 10908
rect 5390 10848 5454 10852
rect 5470 10908 5534 10912
rect 5470 10852 5474 10908
rect 5474 10852 5530 10908
rect 5530 10852 5534 10908
rect 5470 10848 5534 10852
rect 5550 10908 5614 10912
rect 5550 10852 5554 10908
rect 5554 10852 5610 10908
rect 5610 10852 5614 10908
rect 5550 10848 5614 10852
rect 5630 10908 5694 10912
rect 5630 10852 5634 10908
rect 5634 10852 5690 10908
rect 5690 10852 5694 10908
rect 5630 10848 5694 10852
rect 9829 10908 9893 10912
rect 9829 10852 9833 10908
rect 9833 10852 9889 10908
rect 9889 10852 9893 10908
rect 9829 10848 9893 10852
rect 9909 10908 9973 10912
rect 9909 10852 9913 10908
rect 9913 10852 9969 10908
rect 9969 10852 9973 10908
rect 9909 10848 9973 10852
rect 9989 10908 10053 10912
rect 9989 10852 9993 10908
rect 9993 10852 10049 10908
rect 10049 10852 10053 10908
rect 9989 10848 10053 10852
rect 10069 10908 10133 10912
rect 10069 10852 10073 10908
rect 10073 10852 10129 10908
rect 10129 10852 10133 10908
rect 10069 10848 10133 10852
rect 14268 10908 14332 10912
rect 14268 10852 14272 10908
rect 14272 10852 14328 10908
rect 14328 10852 14332 10908
rect 14268 10848 14332 10852
rect 14348 10908 14412 10912
rect 14348 10852 14352 10908
rect 14352 10852 14408 10908
rect 14408 10852 14412 10908
rect 14348 10848 14412 10852
rect 14428 10908 14492 10912
rect 14428 10852 14432 10908
rect 14432 10852 14488 10908
rect 14488 10852 14492 10908
rect 14428 10848 14492 10852
rect 14508 10908 14572 10912
rect 14508 10852 14512 10908
rect 14512 10852 14568 10908
rect 14568 10852 14572 10908
rect 14508 10848 14572 10852
rect 18707 10908 18771 10912
rect 18707 10852 18711 10908
rect 18711 10852 18767 10908
rect 18767 10852 18771 10908
rect 18707 10848 18771 10852
rect 18787 10908 18851 10912
rect 18787 10852 18791 10908
rect 18791 10852 18847 10908
rect 18847 10852 18851 10908
rect 18787 10848 18851 10852
rect 18867 10908 18931 10912
rect 18867 10852 18871 10908
rect 18871 10852 18927 10908
rect 18927 10852 18931 10908
rect 18867 10848 18931 10852
rect 18947 10908 19011 10912
rect 18947 10852 18951 10908
rect 18951 10852 19007 10908
rect 19007 10852 19011 10908
rect 18947 10848 19011 10852
rect 3171 10364 3235 10368
rect 3171 10308 3175 10364
rect 3175 10308 3231 10364
rect 3231 10308 3235 10364
rect 3171 10304 3235 10308
rect 3251 10364 3315 10368
rect 3251 10308 3255 10364
rect 3255 10308 3311 10364
rect 3311 10308 3315 10364
rect 3251 10304 3315 10308
rect 3331 10364 3395 10368
rect 3331 10308 3335 10364
rect 3335 10308 3391 10364
rect 3391 10308 3395 10364
rect 3331 10304 3395 10308
rect 3411 10364 3475 10368
rect 3411 10308 3415 10364
rect 3415 10308 3471 10364
rect 3471 10308 3475 10364
rect 3411 10304 3475 10308
rect 7610 10364 7674 10368
rect 7610 10308 7614 10364
rect 7614 10308 7670 10364
rect 7670 10308 7674 10364
rect 7610 10304 7674 10308
rect 7690 10364 7754 10368
rect 7690 10308 7694 10364
rect 7694 10308 7750 10364
rect 7750 10308 7754 10364
rect 7690 10304 7754 10308
rect 7770 10364 7834 10368
rect 7770 10308 7774 10364
rect 7774 10308 7830 10364
rect 7830 10308 7834 10364
rect 7770 10304 7834 10308
rect 7850 10364 7914 10368
rect 7850 10308 7854 10364
rect 7854 10308 7910 10364
rect 7910 10308 7914 10364
rect 7850 10304 7914 10308
rect 12049 10364 12113 10368
rect 12049 10308 12053 10364
rect 12053 10308 12109 10364
rect 12109 10308 12113 10364
rect 12049 10304 12113 10308
rect 12129 10364 12193 10368
rect 12129 10308 12133 10364
rect 12133 10308 12189 10364
rect 12189 10308 12193 10364
rect 12129 10304 12193 10308
rect 12209 10364 12273 10368
rect 12209 10308 12213 10364
rect 12213 10308 12269 10364
rect 12269 10308 12273 10364
rect 12209 10304 12273 10308
rect 12289 10364 12353 10368
rect 12289 10308 12293 10364
rect 12293 10308 12349 10364
rect 12349 10308 12353 10364
rect 12289 10304 12353 10308
rect 16488 10364 16552 10368
rect 16488 10308 16492 10364
rect 16492 10308 16548 10364
rect 16548 10308 16552 10364
rect 16488 10304 16552 10308
rect 16568 10364 16632 10368
rect 16568 10308 16572 10364
rect 16572 10308 16628 10364
rect 16628 10308 16632 10364
rect 16568 10304 16632 10308
rect 16648 10364 16712 10368
rect 16648 10308 16652 10364
rect 16652 10308 16708 10364
rect 16708 10308 16712 10364
rect 16648 10304 16712 10308
rect 16728 10364 16792 10368
rect 16728 10308 16732 10364
rect 16732 10308 16788 10364
rect 16788 10308 16792 10364
rect 16728 10304 16792 10308
rect 5390 9820 5454 9824
rect 5390 9764 5394 9820
rect 5394 9764 5450 9820
rect 5450 9764 5454 9820
rect 5390 9760 5454 9764
rect 5470 9820 5534 9824
rect 5470 9764 5474 9820
rect 5474 9764 5530 9820
rect 5530 9764 5534 9820
rect 5470 9760 5534 9764
rect 5550 9820 5614 9824
rect 5550 9764 5554 9820
rect 5554 9764 5610 9820
rect 5610 9764 5614 9820
rect 5550 9760 5614 9764
rect 5630 9820 5694 9824
rect 5630 9764 5634 9820
rect 5634 9764 5690 9820
rect 5690 9764 5694 9820
rect 5630 9760 5694 9764
rect 9829 9820 9893 9824
rect 9829 9764 9833 9820
rect 9833 9764 9889 9820
rect 9889 9764 9893 9820
rect 9829 9760 9893 9764
rect 9909 9820 9973 9824
rect 9909 9764 9913 9820
rect 9913 9764 9969 9820
rect 9969 9764 9973 9820
rect 9909 9760 9973 9764
rect 9989 9820 10053 9824
rect 9989 9764 9993 9820
rect 9993 9764 10049 9820
rect 10049 9764 10053 9820
rect 9989 9760 10053 9764
rect 10069 9820 10133 9824
rect 10069 9764 10073 9820
rect 10073 9764 10129 9820
rect 10129 9764 10133 9820
rect 10069 9760 10133 9764
rect 14268 9820 14332 9824
rect 14268 9764 14272 9820
rect 14272 9764 14328 9820
rect 14328 9764 14332 9820
rect 14268 9760 14332 9764
rect 14348 9820 14412 9824
rect 14348 9764 14352 9820
rect 14352 9764 14408 9820
rect 14408 9764 14412 9820
rect 14348 9760 14412 9764
rect 14428 9820 14492 9824
rect 14428 9764 14432 9820
rect 14432 9764 14488 9820
rect 14488 9764 14492 9820
rect 14428 9760 14492 9764
rect 14508 9820 14572 9824
rect 14508 9764 14512 9820
rect 14512 9764 14568 9820
rect 14568 9764 14572 9820
rect 14508 9760 14572 9764
rect 18707 9820 18771 9824
rect 18707 9764 18711 9820
rect 18711 9764 18767 9820
rect 18767 9764 18771 9820
rect 18707 9760 18771 9764
rect 18787 9820 18851 9824
rect 18787 9764 18791 9820
rect 18791 9764 18847 9820
rect 18847 9764 18851 9820
rect 18787 9760 18851 9764
rect 18867 9820 18931 9824
rect 18867 9764 18871 9820
rect 18871 9764 18927 9820
rect 18927 9764 18931 9820
rect 18867 9760 18931 9764
rect 18947 9820 19011 9824
rect 18947 9764 18951 9820
rect 18951 9764 19007 9820
rect 19007 9764 19011 9820
rect 18947 9760 19011 9764
rect 3171 9276 3235 9280
rect 3171 9220 3175 9276
rect 3175 9220 3231 9276
rect 3231 9220 3235 9276
rect 3171 9216 3235 9220
rect 3251 9276 3315 9280
rect 3251 9220 3255 9276
rect 3255 9220 3311 9276
rect 3311 9220 3315 9276
rect 3251 9216 3315 9220
rect 3331 9276 3395 9280
rect 3331 9220 3335 9276
rect 3335 9220 3391 9276
rect 3391 9220 3395 9276
rect 3331 9216 3395 9220
rect 3411 9276 3475 9280
rect 3411 9220 3415 9276
rect 3415 9220 3471 9276
rect 3471 9220 3475 9276
rect 3411 9216 3475 9220
rect 7610 9276 7674 9280
rect 7610 9220 7614 9276
rect 7614 9220 7670 9276
rect 7670 9220 7674 9276
rect 7610 9216 7674 9220
rect 7690 9276 7754 9280
rect 7690 9220 7694 9276
rect 7694 9220 7750 9276
rect 7750 9220 7754 9276
rect 7690 9216 7754 9220
rect 7770 9276 7834 9280
rect 7770 9220 7774 9276
rect 7774 9220 7830 9276
rect 7830 9220 7834 9276
rect 7770 9216 7834 9220
rect 7850 9276 7914 9280
rect 7850 9220 7854 9276
rect 7854 9220 7910 9276
rect 7910 9220 7914 9276
rect 7850 9216 7914 9220
rect 12049 9276 12113 9280
rect 12049 9220 12053 9276
rect 12053 9220 12109 9276
rect 12109 9220 12113 9276
rect 12049 9216 12113 9220
rect 12129 9276 12193 9280
rect 12129 9220 12133 9276
rect 12133 9220 12189 9276
rect 12189 9220 12193 9276
rect 12129 9216 12193 9220
rect 12209 9276 12273 9280
rect 12209 9220 12213 9276
rect 12213 9220 12269 9276
rect 12269 9220 12273 9276
rect 12209 9216 12273 9220
rect 12289 9276 12353 9280
rect 12289 9220 12293 9276
rect 12293 9220 12349 9276
rect 12349 9220 12353 9276
rect 12289 9216 12353 9220
rect 16488 9276 16552 9280
rect 16488 9220 16492 9276
rect 16492 9220 16548 9276
rect 16548 9220 16552 9276
rect 16488 9216 16552 9220
rect 16568 9276 16632 9280
rect 16568 9220 16572 9276
rect 16572 9220 16628 9276
rect 16628 9220 16632 9276
rect 16568 9216 16632 9220
rect 16648 9276 16712 9280
rect 16648 9220 16652 9276
rect 16652 9220 16708 9276
rect 16708 9220 16712 9276
rect 16648 9216 16712 9220
rect 16728 9276 16792 9280
rect 16728 9220 16732 9276
rect 16732 9220 16788 9276
rect 16788 9220 16792 9276
rect 16728 9216 16792 9220
rect 5390 8732 5454 8736
rect 5390 8676 5394 8732
rect 5394 8676 5450 8732
rect 5450 8676 5454 8732
rect 5390 8672 5454 8676
rect 5470 8732 5534 8736
rect 5470 8676 5474 8732
rect 5474 8676 5530 8732
rect 5530 8676 5534 8732
rect 5470 8672 5534 8676
rect 5550 8732 5614 8736
rect 5550 8676 5554 8732
rect 5554 8676 5610 8732
rect 5610 8676 5614 8732
rect 5550 8672 5614 8676
rect 5630 8732 5694 8736
rect 5630 8676 5634 8732
rect 5634 8676 5690 8732
rect 5690 8676 5694 8732
rect 5630 8672 5694 8676
rect 9829 8732 9893 8736
rect 9829 8676 9833 8732
rect 9833 8676 9889 8732
rect 9889 8676 9893 8732
rect 9829 8672 9893 8676
rect 9909 8732 9973 8736
rect 9909 8676 9913 8732
rect 9913 8676 9969 8732
rect 9969 8676 9973 8732
rect 9909 8672 9973 8676
rect 9989 8732 10053 8736
rect 9989 8676 9993 8732
rect 9993 8676 10049 8732
rect 10049 8676 10053 8732
rect 9989 8672 10053 8676
rect 10069 8732 10133 8736
rect 10069 8676 10073 8732
rect 10073 8676 10129 8732
rect 10129 8676 10133 8732
rect 10069 8672 10133 8676
rect 14268 8732 14332 8736
rect 14268 8676 14272 8732
rect 14272 8676 14328 8732
rect 14328 8676 14332 8732
rect 14268 8672 14332 8676
rect 14348 8732 14412 8736
rect 14348 8676 14352 8732
rect 14352 8676 14408 8732
rect 14408 8676 14412 8732
rect 14348 8672 14412 8676
rect 14428 8732 14492 8736
rect 14428 8676 14432 8732
rect 14432 8676 14488 8732
rect 14488 8676 14492 8732
rect 14428 8672 14492 8676
rect 14508 8732 14572 8736
rect 14508 8676 14512 8732
rect 14512 8676 14568 8732
rect 14568 8676 14572 8732
rect 14508 8672 14572 8676
rect 18707 8732 18771 8736
rect 18707 8676 18711 8732
rect 18711 8676 18767 8732
rect 18767 8676 18771 8732
rect 18707 8672 18771 8676
rect 18787 8732 18851 8736
rect 18787 8676 18791 8732
rect 18791 8676 18847 8732
rect 18847 8676 18851 8732
rect 18787 8672 18851 8676
rect 18867 8732 18931 8736
rect 18867 8676 18871 8732
rect 18871 8676 18927 8732
rect 18927 8676 18931 8732
rect 18867 8672 18931 8676
rect 18947 8732 19011 8736
rect 18947 8676 18951 8732
rect 18951 8676 19007 8732
rect 19007 8676 19011 8732
rect 18947 8672 19011 8676
rect 3171 8188 3235 8192
rect 3171 8132 3175 8188
rect 3175 8132 3231 8188
rect 3231 8132 3235 8188
rect 3171 8128 3235 8132
rect 3251 8188 3315 8192
rect 3251 8132 3255 8188
rect 3255 8132 3311 8188
rect 3311 8132 3315 8188
rect 3251 8128 3315 8132
rect 3331 8188 3395 8192
rect 3331 8132 3335 8188
rect 3335 8132 3391 8188
rect 3391 8132 3395 8188
rect 3331 8128 3395 8132
rect 3411 8188 3475 8192
rect 3411 8132 3415 8188
rect 3415 8132 3471 8188
rect 3471 8132 3475 8188
rect 3411 8128 3475 8132
rect 7610 8188 7674 8192
rect 7610 8132 7614 8188
rect 7614 8132 7670 8188
rect 7670 8132 7674 8188
rect 7610 8128 7674 8132
rect 7690 8188 7754 8192
rect 7690 8132 7694 8188
rect 7694 8132 7750 8188
rect 7750 8132 7754 8188
rect 7690 8128 7754 8132
rect 7770 8188 7834 8192
rect 7770 8132 7774 8188
rect 7774 8132 7830 8188
rect 7830 8132 7834 8188
rect 7770 8128 7834 8132
rect 7850 8188 7914 8192
rect 7850 8132 7854 8188
rect 7854 8132 7910 8188
rect 7910 8132 7914 8188
rect 7850 8128 7914 8132
rect 12049 8188 12113 8192
rect 12049 8132 12053 8188
rect 12053 8132 12109 8188
rect 12109 8132 12113 8188
rect 12049 8128 12113 8132
rect 12129 8188 12193 8192
rect 12129 8132 12133 8188
rect 12133 8132 12189 8188
rect 12189 8132 12193 8188
rect 12129 8128 12193 8132
rect 12209 8188 12273 8192
rect 12209 8132 12213 8188
rect 12213 8132 12269 8188
rect 12269 8132 12273 8188
rect 12209 8128 12273 8132
rect 12289 8188 12353 8192
rect 12289 8132 12293 8188
rect 12293 8132 12349 8188
rect 12349 8132 12353 8188
rect 12289 8128 12353 8132
rect 16488 8188 16552 8192
rect 16488 8132 16492 8188
rect 16492 8132 16548 8188
rect 16548 8132 16552 8188
rect 16488 8128 16552 8132
rect 16568 8188 16632 8192
rect 16568 8132 16572 8188
rect 16572 8132 16628 8188
rect 16628 8132 16632 8188
rect 16568 8128 16632 8132
rect 16648 8188 16712 8192
rect 16648 8132 16652 8188
rect 16652 8132 16708 8188
rect 16708 8132 16712 8188
rect 16648 8128 16712 8132
rect 16728 8188 16792 8192
rect 16728 8132 16732 8188
rect 16732 8132 16788 8188
rect 16788 8132 16792 8188
rect 16728 8128 16792 8132
rect 5390 7644 5454 7648
rect 5390 7588 5394 7644
rect 5394 7588 5450 7644
rect 5450 7588 5454 7644
rect 5390 7584 5454 7588
rect 5470 7644 5534 7648
rect 5470 7588 5474 7644
rect 5474 7588 5530 7644
rect 5530 7588 5534 7644
rect 5470 7584 5534 7588
rect 5550 7644 5614 7648
rect 5550 7588 5554 7644
rect 5554 7588 5610 7644
rect 5610 7588 5614 7644
rect 5550 7584 5614 7588
rect 5630 7644 5694 7648
rect 5630 7588 5634 7644
rect 5634 7588 5690 7644
rect 5690 7588 5694 7644
rect 5630 7584 5694 7588
rect 9829 7644 9893 7648
rect 9829 7588 9833 7644
rect 9833 7588 9889 7644
rect 9889 7588 9893 7644
rect 9829 7584 9893 7588
rect 9909 7644 9973 7648
rect 9909 7588 9913 7644
rect 9913 7588 9969 7644
rect 9969 7588 9973 7644
rect 9909 7584 9973 7588
rect 9989 7644 10053 7648
rect 9989 7588 9993 7644
rect 9993 7588 10049 7644
rect 10049 7588 10053 7644
rect 9989 7584 10053 7588
rect 10069 7644 10133 7648
rect 10069 7588 10073 7644
rect 10073 7588 10129 7644
rect 10129 7588 10133 7644
rect 10069 7584 10133 7588
rect 14268 7644 14332 7648
rect 14268 7588 14272 7644
rect 14272 7588 14328 7644
rect 14328 7588 14332 7644
rect 14268 7584 14332 7588
rect 14348 7644 14412 7648
rect 14348 7588 14352 7644
rect 14352 7588 14408 7644
rect 14408 7588 14412 7644
rect 14348 7584 14412 7588
rect 14428 7644 14492 7648
rect 14428 7588 14432 7644
rect 14432 7588 14488 7644
rect 14488 7588 14492 7644
rect 14428 7584 14492 7588
rect 14508 7644 14572 7648
rect 14508 7588 14512 7644
rect 14512 7588 14568 7644
rect 14568 7588 14572 7644
rect 14508 7584 14572 7588
rect 18707 7644 18771 7648
rect 18707 7588 18711 7644
rect 18711 7588 18767 7644
rect 18767 7588 18771 7644
rect 18707 7584 18771 7588
rect 18787 7644 18851 7648
rect 18787 7588 18791 7644
rect 18791 7588 18847 7644
rect 18847 7588 18851 7644
rect 18787 7584 18851 7588
rect 18867 7644 18931 7648
rect 18867 7588 18871 7644
rect 18871 7588 18927 7644
rect 18927 7588 18931 7644
rect 18867 7584 18931 7588
rect 18947 7644 19011 7648
rect 18947 7588 18951 7644
rect 18951 7588 19007 7644
rect 19007 7588 19011 7644
rect 18947 7584 19011 7588
rect 3171 7100 3235 7104
rect 3171 7044 3175 7100
rect 3175 7044 3231 7100
rect 3231 7044 3235 7100
rect 3171 7040 3235 7044
rect 3251 7100 3315 7104
rect 3251 7044 3255 7100
rect 3255 7044 3311 7100
rect 3311 7044 3315 7100
rect 3251 7040 3315 7044
rect 3331 7100 3395 7104
rect 3331 7044 3335 7100
rect 3335 7044 3391 7100
rect 3391 7044 3395 7100
rect 3331 7040 3395 7044
rect 3411 7100 3475 7104
rect 3411 7044 3415 7100
rect 3415 7044 3471 7100
rect 3471 7044 3475 7100
rect 3411 7040 3475 7044
rect 7610 7100 7674 7104
rect 7610 7044 7614 7100
rect 7614 7044 7670 7100
rect 7670 7044 7674 7100
rect 7610 7040 7674 7044
rect 7690 7100 7754 7104
rect 7690 7044 7694 7100
rect 7694 7044 7750 7100
rect 7750 7044 7754 7100
rect 7690 7040 7754 7044
rect 7770 7100 7834 7104
rect 7770 7044 7774 7100
rect 7774 7044 7830 7100
rect 7830 7044 7834 7100
rect 7770 7040 7834 7044
rect 7850 7100 7914 7104
rect 7850 7044 7854 7100
rect 7854 7044 7910 7100
rect 7910 7044 7914 7100
rect 7850 7040 7914 7044
rect 12049 7100 12113 7104
rect 12049 7044 12053 7100
rect 12053 7044 12109 7100
rect 12109 7044 12113 7100
rect 12049 7040 12113 7044
rect 12129 7100 12193 7104
rect 12129 7044 12133 7100
rect 12133 7044 12189 7100
rect 12189 7044 12193 7100
rect 12129 7040 12193 7044
rect 12209 7100 12273 7104
rect 12209 7044 12213 7100
rect 12213 7044 12269 7100
rect 12269 7044 12273 7100
rect 12209 7040 12273 7044
rect 12289 7100 12353 7104
rect 12289 7044 12293 7100
rect 12293 7044 12349 7100
rect 12349 7044 12353 7100
rect 12289 7040 12353 7044
rect 16488 7100 16552 7104
rect 16488 7044 16492 7100
rect 16492 7044 16548 7100
rect 16548 7044 16552 7100
rect 16488 7040 16552 7044
rect 16568 7100 16632 7104
rect 16568 7044 16572 7100
rect 16572 7044 16628 7100
rect 16628 7044 16632 7100
rect 16568 7040 16632 7044
rect 16648 7100 16712 7104
rect 16648 7044 16652 7100
rect 16652 7044 16708 7100
rect 16708 7044 16712 7100
rect 16648 7040 16712 7044
rect 16728 7100 16792 7104
rect 16728 7044 16732 7100
rect 16732 7044 16788 7100
rect 16788 7044 16792 7100
rect 16728 7040 16792 7044
rect 5390 6556 5454 6560
rect 5390 6500 5394 6556
rect 5394 6500 5450 6556
rect 5450 6500 5454 6556
rect 5390 6496 5454 6500
rect 5470 6556 5534 6560
rect 5470 6500 5474 6556
rect 5474 6500 5530 6556
rect 5530 6500 5534 6556
rect 5470 6496 5534 6500
rect 5550 6556 5614 6560
rect 5550 6500 5554 6556
rect 5554 6500 5610 6556
rect 5610 6500 5614 6556
rect 5550 6496 5614 6500
rect 5630 6556 5694 6560
rect 5630 6500 5634 6556
rect 5634 6500 5690 6556
rect 5690 6500 5694 6556
rect 5630 6496 5694 6500
rect 9829 6556 9893 6560
rect 9829 6500 9833 6556
rect 9833 6500 9889 6556
rect 9889 6500 9893 6556
rect 9829 6496 9893 6500
rect 9909 6556 9973 6560
rect 9909 6500 9913 6556
rect 9913 6500 9969 6556
rect 9969 6500 9973 6556
rect 9909 6496 9973 6500
rect 9989 6556 10053 6560
rect 9989 6500 9993 6556
rect 9993 6500 10049 6556
rect 10049 6500 10053 6556
rect 9989 6496 10053 6500
rect 10069 6556 10133 6560
rect 10069 6500 10073 6556
rect 10073 6500 10129 6556
rect 10129 6500 10133 6556
rect 10069 6496 10133 6500
rect 14268 6556 14332 6560
rect 14268 6500 14272 6556
rect 14272 6500 14328 6556
rect 14328 6500 14332 6556
rect 14268 6496 14332 6500
rect 14348 6556 14412 6560
rect 14348 6500 14352 6556
rect 14352 6500 14408 6556
rect 14408 6500 14412 6556
rect 14348 6496 14412 6500
rect 14428 6556 14492 6560
rect 14428 6500 14432 6556
rect 14432 6500 14488 6556
rect 14488 6500 14492 6556
rect 14428 6496 14492 6500
rect 14508 6556 14572 6560
rect 14508 6500 14512 6556
rect 14512 6500 14568 6556
rect 14568 6500 14572 6556
rect 14508 6496 14572 6500
rect 18707 6556 18771 6560
rect 18707 6500 18711 6556
rect 18711 6500 18767 6556
rect 18767 6500 18771 6556
rect 18707 6496 18771 6500
rect 18787 6556 18851 6560
rect 18787 6500 18791 6556
rect 18791 6500 18847 6556
rect 18847 6500 18851 6556
rect 18787 6496 18851 6500
rect 18867 6556 18931 6560
rect 18867 6500 18871 6556
rect 18871 6500 18927 6556
rect 18927 6500 18931 6556
rect 18867 6496 18931 6500
rect 18947 6556 19011 6560
rect 18947 6500 18951 6556
rect 18951 6500 19007 6556
rect 19007 6500 19011 6556
rect 18947 6496 19011 6500
rect 3171 6012 3235 6016
rect 3171 5956 3175 6012
rect 3175 5956 3231 6012
rect 3231 5956 3235 6012
rect 3171 5952 3235 5956
rect 3251 6012 3315 6016
rect 3251 5956 3255 6012
rect 3255 5956 3311 6012
rect 3311 5956 3315 6012
rect 3251 5952 3315 5956
rect 3331 6012 3395 6016
rect 3331 5956 3335 6012
rect 3335 5956 3391 6012
rect 3391 5956 3395 6012
rect 3331 5952 3395 5956
rect 3411 6012 3475 6016
rect 3411 5956 3415 6012
rect 3415 5956 3471 6012
rect 3471 5956 3475 6012
rect 3411 5952 3475 5956
rect 7610 6012 7674 6016
rect 7610 5956 7614 6012
rect 7614 5956 7670 6012
rect 7670 5956 7674 6012
rect 7610 5952 7674 5956
rect 7690 6012 7754 6016
rect 7690 5956 7694 6012
rect 7694 5956 7750 6012
rect 7750 5956 7754 6012
rect 7690 5952 7754 5956
rect 7770 6012 7834 6016
rect 7770 5956 7774 6012
rect 7774 5956 7830 6012
rect 7830 5956 7834 6012
rect 7770 5952 7834 5956
rect 7850 6012 7914 6016
rect 7850 5956 7854 6012
rect 7854 5956 7910 6012
rect 7910 5956 7914 6012
rect 7850 5952 7914 5956
rect 12049 6012 12113 6016
rect 12049 5956 12053 6012
rect 12053 5956 12109 6012
rect 12109 5956 12113 6012
rect 12049 5952 12113 5956
rect 12129 6012 12193 6016
rect 12129 5956 12133 6012
rect 12133 5956 12189 6012
rect 12189 5956 12193 6012
rect 12129 5952 12193 5956
rect 12209 6012 12273 6016
rect 12209 5956 12213 6012
rect 12213 5956 12269 6012
rect 12269 5956 12273 6012
rect 12209 5952 12273 5956
rect 12289 6012 12353 6016
rect 12289 5956 12293 6012
rect 12293 5956 12349 6012
rect 12349 5956 12353 6012
rect 12289 5952 12353 5956
rect 16488 6012 16552 6016
rect 16488 5956 16492 6012
rect 16492 5956 16548 6012
rect 16548 5956 16552 6012
rect 16488 5952 16552 5956
rect 16568 6012 16632 6016
rect 16568 5956 16572 6012
rect 16572 5956 16628 6012
rect 16628 5956 16632 6012
rect 16568 5952 16632 5956
rect 16648 6012 16712 6016
rect 16648 5956 16652 6012
rect 16652 5956 16708 6012
rect 16708 5956 16712 6012
rect 16648 5952 16712 5956
rect 16728 6012 16792 6016
rect 16728 5956 16732 6012
rect 16732 5956 16788 6012
rect 16788 5956 16792 6012
rect 16728 5952 16792 5956
rect 5390 5468 5454 5472
rect 5390 5412 5394 5468
rect 5394 5412 5450 5468
rect 5450 5412 5454 5468
rect 5390 5408 5454 5412
rect 5470 5468 5534 5472
rect 5470 5412 5474 5468
rect 5474 5412 5530 5468
rect 5530 5412 5534 5468
rect 5470 5408 5534 5412
rect 5550 5468 5614 5472
rect 5550 5412 5554 5468
rect 5554 5412 5610 5468
rect 5610 5412 5614 5468
rect 5550 5408 5614 5412
rect 5630 5468 5694 5472
rect 5630 5412 5634 5468
rect 5634 5412 5690 5468
rect 5690 5412 5694 5468
rect 5630 5408 5694 5412
rect 9829 5468 9893 5472
rect 9829 5412 9833 5468
rect 9833 5412 9889 5468
rect 9889 5412 9893 5468
rect 9829 5408 9893 5412
rect 9909 5468 9973 5472
rect 9909 5412 9913 5468
rect 9913 5412 9969 5468
rect 9969 5412 9973 5468
rect 9909 5408 9973 5412
rect 9989 5468 10053 5472
rect 9989 5412 9993 5468
rect 9993 5412 10049 5468
rect 10049 5412 10053 5468
rect 9989 5408 10053 5412
rect 10069 5468 10133 5472
rect 10069 5412 10073 5468
rect 10073 5412 10129 5468
rect 10129 5412 10133 5468
rect 10069 5408 10133 5412
rect 14268 5468 14332 5472
rect 14268 5412 14272 5468
rect 14272 5412 14328 5468
rect 14328 5412 14332 5468
rect 14268 5408 14332 5412
rect 14348 5468 14412 5472
rect 14348 5412 14352 5468
rect 14352 5412 14408 5468
rect 14408 5412 14412 5468
rect 14348 5408 14412 5412
rect 14428 5468 14492 5472
rect 14428 5412 14432 5468
rect 14432 5412 14488 5468
rect 14488 5412 14492 5468
rect 14428 5408 14492 5412
rect 14508 5468 14572 5472
rect 14508 5412 14512 5468
rect 14512 5412 14568 5468
rect 14568 5412 14572 5468
rect 14508 5408 14572 5412
rect 18707 5468 18771 5472
rect 18707 5412 18711 5468
rect 18711 5412 18767 5468
rect 18767 5412 18771 5468
rect 18707 5408 18771 5412
rect 18787 5468 18851 5472
rect 18787 5412 18791 5468
rect 18791 5412 18847 5468
rect 18847 5412 18851 5468
rect 18787 5408 18851 5412
rect 18867 5468 18931 5472
rect 18867 5412 18871 5468
rect 18871 5412 18927 5468
rect 18927 5412 18931 5468
rect 18867 5408 18931 5412
rect 18947 5468 19011 5472
rect 18947 5412 18951 5468
rect 18951 5412 19007 5468
rect 19007 5412 19011 5468
rect 18947 5408 19011 5412
rect 3171 4924 3235 4928
rect 3171 4868 3175 4924
rect 3175 4868 3231 4924
rect 3231 4868 3235 4924
rect 3171 4864 3235 4868
rect 3251 4924 3315 4928
rect 3251 4868 3255 4924
rect 3255 4868 3311 4924
rect 3311 4868 3315 4924
rect 3251 4864 3315 4868
rect 3331 4924 3395 4928
rect 3331 4868 3335 4924
rect 3335 4868 3391 4924
rect 3391 4868 3395 4924
rect 3331 4864 3395 4868
rect 3411 4924 3475 4928
rect 3411 4868 3415 4924
rect 3415 4868 3471 4924
rect 3471 4868 3475 4924
rect 3411 4864 3475 4868
rect 7610 4924 7674 4928
rect 7610 4868 7614 4924
rect 7614 4868 7670 4924
rect 7670 4868 7674 4924
rect 7610 4864 7674 4868
rect 7690 4924 7754 4928
rect 7690 4868 7694 4924
rect 7694 4868 7750 4924
rect 7750 4868 7754 4924
rect 7690 4864 7754 4868
rect 7770 4924 7834 4928
rect 7770 4868 7774 4924
rect 7774 4868 7830 4924
rect 7830 4868 7834 4924
rect 7770 4864 7834 4868
rect 7850 4924 7914 4928
rect 7850 4868 7854 4924
rect 7854 4868 7910 4924
rect 7910 4868 7914 4924
rect 7850 4864 7914 4868
rect 12049 4924 12113 4928
rect 12049 4868 12053 4924
rect 12053 4868 12109 4924
rect 12109 4868 12113 4924
rect 12049 4864 12113 4868
rect 12129 4924 12193 4928
rect 12129 4868 12133 4924
rect 12133 4868 12189 4924
rect 12189 4868 12193 4924
rect 12129 4864 12193 4868
rect 12209 4924 12273 4928
rect 12209 4868 12213 4924
rect 12213 4868 12269 4924
rect 12269 4868 12273 4924
rect 12209 4864 12273 4868
rect 12289 4924 12353 4928
rect 12289 4868 12293 4924
rect 12293 4868 12349 4924
rect 12349 4868 12353 4924
rect 12289 4864 12353 4868
rect 16488 4924 16552 4928
rect 16488 4868 16492 4924
rect 16492 4868 16548 4924
rect 16548 4868 16552 4924
rect 16488 4864 16552 4868
rect 16568 4924 16632 4928
rect 16568 4868 16572 4924
rect 16572 4868 16628 4924
rect 16628 4868 16632 4924
rect 16568 4864 16632 4868
rect 16648 4924 16712 4928
rect 16648 4868 16652 4924
rect 16652 4868 16708 4924
rect 16708 4868 16712 4924
rect 16648 4864 16712 4868
rect 16728 4924 16792 4928
rect 16728 4868 16732 4924
rect 16732 4868 16788 4924
rect 16788 4868 16792 4924
rect 16728 4864 16792 4868
rect 5390 4380 5454 4384
rect 5390 4324 5394 4380
rect 5394 4324 5450 4380
rect 5450 4324 5454 4380
rect 5390 4320 5454 4324
rect 5470 4380 5534 4384
rect 5470 4324 5474 4380
rect 5474 4324 5530 4380
rect 5530 4324 5534 4380
rect 5470 4320 5534 4324
rect 5550 4380 5614 4384
rect 5550 4324 5554 4380
rect 5554 4324 5610 4380
rect 5610 4324 5614 4380
rect 5550 4320 5614 4324
rect 5630 4380 5694 4384
rect 5630 4324 5634 4380
rect 5634 4324 5690 4380
rect 5690 4324 5694 4380
rect 5630 4320 5694 4324
rect 9829 4380 9893 4384
rect 9829 4324 9833 4380
rect 9833 4324 9889 4380
rect 9889 4324 9893 4380
rect 9829 4320 9893 4324
rect 9909 4380 9973 4384
rect 9909 4324 9913 4380
rect 9913 4324 9969 4380
rect 9969 4324 9973 4380
rect 9909 4320 9973 4324
rect 9989 4380 10053 4384
rect 9989 4324 9993 4380
rect 9993 4324 10049 4380
rect 10049 4324 10053 4380
rect 9989 4320 10053 4324
rect 10069 4380 10133 4384
rect 10069 4324 10073 4380
rect 10073 4324 10129 4380
rect 10129 4324 10133 4380
rect 10069 4320 10133 4324
rect 14268 4380 14332 4384
rect 14268 4324 14272 4380
rect 14272 4324 14328 4380
rect 14328 4324 14332 4380
rect 14268 4320 14332 4324
rect 14348 4380 14412 4384
rect 14348 4324 14352 4380
rect 14352 4324 14408 4380
rect 14408 4324 14412 4380
rect 14348 4320 14412 4324
rect 14428 4380 14492 4384
rect 14428 4324 14432 4380
rect 14432 4324 14488 4380
rect 14488 4324 14492 4380
rect 14428 4320 14492 4324
rect 14508 4380 14572 4384
rect 14508 4324 14512 4380
rect 14512 4324 14568 4380
rect 14568 4324 14572 4380
rect 14508 4320 14572 4324
rect 18707 4380 18771 4384
rect 18707 4324 18711 4380
rect 18711 4324 18767 4380
rect 18767 4324 18771 4380
rect 18707 4320 18771 4324
rect 18787 4380 18851 4384
rect 18787 4324 18791 4380
rect 18791 4324 18847 4380
rect 18847 4324 18851 4380
rect 18787 4320 18851 4324
rect 18867 4380 18931 4384
rect 18867 4324 18871 4380
rect 18871 4324 18927 4380
rect 18927 4324 18931 4380
rect 18867 4320 18931 4324
rect 18947 4380 19011 4384
rect 18947 4324 18951 4380
rect 18951 4324 19007 4380
rect 19007 4324 19011 4380
rect 18947 4320 19011 4324
rect 3171 3836 3235 3840
rect 3171 3780 3175 3836
rect 3175 3780 3231 3836
rect 3231 3780 3235 3836
rect 3171 3776 3235 3780
rect 3251 3836 3315 3840
rect 3251 3780 3255 3836
rect 3255 3780 3311 3836
rect 3311 3780 3315 3836
rect 3251 3776 3315 3780
rect 3331 3836 3395 3840
rect 3331 3780 3335 3836
rect 3335 3780 3391 3836
rect 3391 3780 3395 3836
rect 3331 3776 3395 3780
rect 3411 3836 3475 3840
rect 3411 3780 3415 3836
rect 3415 3780 3471 3836
rect 3471 3780 3475 3836
rect 3411 3776 3475 3780
rect 7610 3836 7674 3840
rect 7610 3780 7614 3836
rect 7614 3780 7670 3836
rect 7670 3780 7674 3836
rect 7610 3776 7674 3780
rect 7690 3836 7754 3840
rect 7690 3780 7694 3836
rect 7694 3780 7750 3836
rect 7750 3780 7754 3836
rect 7690 3776 7754 3780
rect 7770 3836 7834 3840
rect 7770 3780 7774 3836
rect 7774 3780 7830 3836
rect 7830 3780 7834 3836
rect 7770 3776 7834 3780
rect 7850 3836 7914 3840
rect 7850 3780 7854 3836
rect 7854 3780 7910 3836
rect 7910 3780 7914 3836
rect 7850 3776 7914 3780
rect 12049 3836 12113 3840
rect 12049 3780 12053 3836
rect 12053 3780 12109 3836
rect 12109 3780 12113 3836
rect 12049 3776 12113 3780
rect 12129 3836 12193 3840
rect 12129 3780 12133 3836
rect 12133 3780 12189 3836
rect 12189 3780 12193 3836
rect 12129 3776 12193 3780
rect 12209 3836 12273 3840
rect 12209 3780 12213 3836
rect 12213 3780 12269 3836
rect 12269 3780 12273 3836
rect 12209 3776 12273 3780
rect 12289 3836 12353 3840
rect 12289 3780 12293 3836
rect 12293 3780 12349 3836
rect 12349 3780 12353 3836
rect 12289 3776 12353 3780
rect 16488 3836 16552 3840
rect 16488 3780 16492 3836
rect 16492 3780 16548 3836
rect 16548 3780 16552 3836
rect 16488 3776 16552 3780
rect 16568 3836 16632 3840
rect 16568 3780 16572 3836
rect 16572 3780 16628 3836
rect 16628 3780 16632 3836
rect 16568 3776 16632 3780
rect 16648 3836 16712 3840
rect 16648 3780 16652 3836
rect 16652 3780 16708 3836
rect 16708 3780 16712 3836
rect 16648 3776 16712 3780
rect 16728 3836 16792 3840
rect 16728 3780 16732 3836
rect 16732 3780 16788 3836
rect 16788 3780 16792 3836
rect 16728 3776 16792 3780
rect 5390 3292 5454 3296
rect 5390 3236 5394 3292
rect 5394 3236 5450 3292
rect 5450 3236 5454 3292
rect 5390 3232 5454 3236
rect 5470 3292 5534 3296
rect 5470 3236 5474 3292
rect 5474 3236 5530 3292
rect 5530 3236 5534 3292
rect 5470 3232 5534 3236
rect 5550 3292 5614 3296
rect 5550 3236 5554 3292
rect 5554 3236 5610 3292
rect 5610 3236 5614 3292
rect 5550 3232 5614 3236
rect 5630 3292 5694 3296
rect 5630 3236 5634 3292
rect 5634 3236 5690 3292
rect 5690 3236 5694 3292
rect 5630 3232 5694 3236
rect 9829 3292 9893 3296
rect 9829 3236 9833 3292
rect 9833 3236 9889 3292
rect 9889 3236 9893 3292
rect 9829 3232 9893 3236
rect 9909 3292 9973 3296
rect 9909 3236 9913 3292
rect 9913 3236 9969 3292
rect 9969 3236 9973 3292
rect 9909 3232 9973 3236
rect 9989 3292 10053 3296
rect 9989 3236 9993 3292
rect 9993 3236 10049 3292
rect 10049 3236 10053 3292
rect 9989 3232 10053 3236
rect 10069 3292 10133 3296
rect 10069 3236 10073 3292
rect 10073 3236 10129 3292
rect 10129 3236 10133 3292
rect 10069 3232 10133 3236
rect 14268 3292 14332 3296
rect 14268 3236 14272 3292
rect 14272 3236 14328 3292
rect 14328 3236 14332 3292
rect 14268 3232 14332 3236
rect 14348 3292 14412 3296
rect 14348 3236 14352 3292
rect 14352 3236 14408 3292
rect 14408 3236 14412 3292
rect 14348 3232 14412 3236
rect 14428 3292 14492 3296
rect 14428 3236 14432 3292
rect 14432 3236 14488 3292
rect 14488 3236 14492 3292
rect 14428 3232 14492 3236
rect 14508 3292 14572 3296
rect 14508 3236 14512 3292
rect 14512 3236 14568 3292
rect 14568 3236 14572 3292
rect 14508 3232 14572 3236
rect 18707 3292 18771 3296
rect 18707 3236 18711 3292
rect 18711 3236 18767 3292
rect 18767 3236 18771 3292
rect 18707 3232 18771 3236
rect 18787 3292 18851 3296
rect 18787 3236 18791 3292
rect 18791 3236 18847 3292
rect 18847 3236 18851 3292
rect 18787 3232 18851 3236
rect 18867 3292 18931 3296
rect 18867 3236 18871 3292
rect 18871 3236 18927 3292
rect 18927 3236 18931 3292
rect 18867 3232 18931 3236
rect 18947 3292 19011 3296
rect 18947 3236 18951 3292
rect 18951 3236 19007 3292
rect 19007 3236 19011 3292
rect 18947 3232 19011 3236
rect 3171 2748 3235 2752
rect 3171 2692 3175 2748
rect 3175 2692 3231 2748
rect 3231 2692 3235 2748
rect 3171 2688 3235 2692
rect 3251 2748 3315 2752
rect 3251 2692 3255 2748
rect 3255 2692 3311 2748
rect 3311 2692 3315 2748
rect 3251 2688 3315 2692
rect 3331 2748 3395 2752
rect 3331 2692 3335 2748
rect 3335 2692 3391 2748
rect 3391 2692 3395 2748
rect 3331 2688 3395 2692
rect 3411 2748 3475 2752
rect 3411 2692 3415 2748
rect 3415 2692 3471 2748
rect 3471 2692 3475 2748
rect 3411 2688 3475 2692
rect 7610 2748 7674 2752
rect 7610 2692 7614 2748
rect 7614 2692 7670 2748
rect 7670 2692 7674 2748
rect 7610 2688 7674 2692
rect 7690 2748 7754 2752
rect 7690 2692 7694 2748
rect 7694 2692 7750 2748
rect 7750 2692 7754 2748
rect 7690 2688 7754 2692
rect 7770 2748 7834 2752
rect 7770 2692 7774 2748
rect 7774 2692 7830 2748
rect 7830 2692 7834 2748
rect 7770 2688 7834 2692
rect 7850 2748 7914 2752
rect 7850 2692 7854 2748
rect 7854 2692 7910 2748
rect 7910 2692 7914 2748
rect 7850 2688 7914 2692
rect 12049 2748 12113 2752
rect 12049 2692 12053 2748
rect 12053 2692 12109 2748
rect 12109 2692 12113 2748
rect 12049 2688 12113 2692
rect 12129 2748 12193 2752
rect 12129 2692 12133 2748
rect 12133 2692 12189 2748
rect 12189 2692 12193 2748
rect 12129 2688 12193 2692
rect 12209 2748 12273 2752
rect 12209 2692 12213 2748
rect 12213 2692 12269 2748
rect 12269 2692 12273 2748
rect 12209 2688 12273 2692
rect 12289 2748 12353 2752
rect 12289 2692 12293 2748
rect 12293 2692 12349 2748
rect 12349 2692 12353 2748
rect 12289 2688 12353 2692
rect 16488 2748 16552 2752
rect 16488 2692 16492 2748
rect 16492 2692 16548 2748
rect 16548 2692 16552 2748
rect 16488 2688 16552 2692
rect 16568 2748 16632 2752
rect 16568 2692 16572 2748
rect 16572 2692 16628 2748
rect 16628 2692 16632 2748
rect 16568 2688 16632 2692
rect 16648 2748 16712 2752
rect 16648 2692 16652 2748
rect 16652 2692 16708 2748
rect 16708 2692 16712 2748
rect 16648 2688 16712 2692
rect 16728 2748 16792 2752
rect 16728 2692 16732 2748
rect 16732 2692 16788 2748
rect 16788 2692 16792 2748
rect 16728 2688 16792 2692
rect 5390 2204 5454 2208
rect 5390 2148 5394 2204
rect 5394 2148 5450 2204
rect 5450 2148 5454 2204
rect 5390 2144 5454 2148
rect 5470 2204 5534 2208
rect 5470 2148 5474 2204
rect 5474 2148 5530 2204
rect 5530 2148 5534 2204
rect 5470 2144 5534 2148
rect 5550 2204 5614 2208
rect 5550 2148 5554 2204
rect 5554 2148 5610 2204
rect 5610 2148 5614 2204
rect 5550 2144 5614 2148
rect 5630 2204 5694 2208
rect 5630 2148 5634 2204
rect 5634 2148 5690 2204
rect 5690 2148 5694 2204
rect 5630 2144 5694 2148
rect 9829 2204 9893 2208
rect 9829 2148 9833 2204
rect 9833 2148 9889 2204
rect 9889 2148 9893 2204
rect 9829 2144 9893 2148
rect 9909 2204 9973 2208
rect 9909 2148 9913 2204
rect 9913 2148 9969 2204
rect 9969 2148 9973 2204
rect 9909 2144 9973 2148
rect 9989 2204 10053 2208
rect 9989 2148 9993 2204
rect 9993 2148 10049 2204
rect 10049 2148 10053 2204
rect 9989 2144 10053 2148
rect 10069 2204 10133 2208
rect 10069 2148 10073 2204
rect 10073 2148 10129 2204
rect 10129 2148 10133 2204
rect 10069 2144 10133 2148
rect 14268 2204 14332 2208
rect 14268 2148 14272 2204
rect 14272 2148 14328 2204
rect 14328 2148 14332 2204
rect 14268 2144 14332 2148
rect 14348 2204 14412 2208
rect 14348 2148 14352 2204
rect 14352 2148 14408 2204
rect 14408 2148 14412 2204
rect 14348 2144 14412 2148
rect 14428 2204 14492 2208
rect 14428 2148 14432 2204
rect 14432 2148 14488 2204
rect 14488 2148 14492 2204
rect 14428 2144 14492 2148
rect 14508 2204 14572 2208
rect 14508 2148 14512 2204
rect 14512 2148 14568 2204
rect 14568 2148 14572 2204
rect 14508 2144 14572 2148
rect 18707 2204 18771 2208
rect 18707 2148 18711 2204
rect 18711 2148 18767 2204
rect 18767 2148 18771 2204
rect 18707 2144 18771 2148
rect 18787 2204 18851 2208
rect 18787 2148 18791 2204
rect 18791 2148 18847 2204
rect 18847 2148 18851 2204
rect 18787 2144 18851 2148
rect 18867 2204 18931 2208
rect 18867 2148 18871 2204
rect 18871 2148 18927 2204
rect 18927 2148 18931 2204
rect 18867 2144 18931 2148
rect 18947 2204 19011 2208
rect 18947 2148 18951 2204
rect 18951 2148 19007 2204
rect 19007 2148 19011 2204
rect 18947 2144 19011 2148
<< metal4 >>
rect 3163 47360 3483 47376
rect 3163 47296 3171 47360
rect 3235 47296 3251 47360
rect 3315 47296 3331 47360
rect 3395 47296 3411 47360
rect 3475 47296 3483 47360
rect 3163 46272 3483 47296
rect 3163 46208 3171 46272
rect 3235 46208 3251 46272
rect 3315 46208 3331 46272
rect 3395 46208 3411 46272
rect 3475 46208 3483 46272
rect 3163 45184 3483 46208
rect 3163 45120 3171 45184
rect 3235 45120 3251 45184
rect 3315 45120 3331 45184
rect 3395 45120 3411 45184
rect 3475 45120 3483 45184
rect 3163 44096 3483 45120
rect 3163 44032 3171 44096
rect 3235 44032 3251 44096
rect 3315 44032 3331 44096
rect 3395 44032 3411 44096
rect 3475 44032 3483 44096
rect 3163 43008 3483 44032
rect 3163 42944 3171 43008
rect 3235 42944 3251 43008
rect 3315 42944 3331 43008
rect 3395 42944 3411 43008
rect 3475 42944 3483 43008
rect 3163 41920 3483 42944
rect 3163 41856 3171 41920
rect 3235 41856 3251 41920
rect 3315 41856 3331 41920
rect 3395 41856 3411 41920
rect 3475 41856 3483 41920
rect 3163 40832 3483 41856
rect 3163 40768 3171 40832
rect 3235 40768 3251 40832
rect 3315 40768 3331 40832
rect 3395 40768 3411 40832
rect 3475 40768 3483 40832
rect 3163 39744 3483 40768
rect 3163 39680 3171 39744
rect 3235 39680 3251 39744
rect 3315 39680 3331 39744
rect 3395 39680 3411 39744
rect 3475 39680 3483 39744
rect 3163 38656 3483 39680
rect 3163 38592 3171 38656
rect 3235 38592 3251 38656
rect 3315 38592 3331 38656
rect 3395 38592 3411 38656
rect 3475 38592 3483 38656
rect 3163 37568 3483 38592
rect 3163 37504 3171 37568
rect 3235 37504 3251 37568
rect 3315 37504 3331 37568
rect 3395 37504 3411 37568
rect 3475 37504 3483 37568
rect 3163 36480 3483 37504
rect 3163 36416 3171 36480
rect 3235 36416 3251 36480
rect 3315 36416 3331 36480
rect 3395 36416 3411 36480
rect 3475 36416 3483 36480
rect 3163 35392 3483 36416
rect 3163 35328 3171 35392
rect 3235 35328 3251 35392
rect 3315 35328 3331 35392
rect 3395 35328 3411 35392
rect 3475 35328 3483 35392
rect 3163 34304 3483 35328
rect 3163 34240 3171 34304
rect 3235 34240 3251 34304
rect 3315 34240 3331 34304
rect 3395 34240 3411 34304
rect 3475 34240 3483 34304
rect 3163 33216 3483 34240
rect 3163 33152 3171 33216
rect 3235 33152 3251 33216
rect 3315 33152 3331 33216
rect 3395 33152 3411 33216
rect 3475 33152 3483 33216
rect 3163 32128 3483 33152
rect 3163 32064 3171 32128
rect 3235 32064 3251 32128
rect 3315 32064 3331 32128
rect 3395 32064 3411 32128
rect 3475 32064 3483 32128
rect 3163 31040 3483 32064
rect 3163 30976 3171 31040
rect 3235 30976 3251 31040
rect 3315 30976 3331 31040
rect 3395 30976 3411 31040
rect 3475 30976 3483 31040
rect 3163 29952 3483 30976
rect 3163 29888 3171 29952
rect 3235 29888 3251 29952
rect 3315 29888 3331 29952
rect 3395 29888 3411 29952
rect 3475 29888 3483 29952
rect 3163 28864 3483 29888
rect 3163 28800 3171 28864
rect 3235 28800 3251 28864
rect 3315 28800 3331 28864
rect 3395 28800 3411 28864
rect 3475 28800 3483 28864
rect 3163 27776 3483 28800
rect 3163 27712 3171 27776
rect 3235 27712 3251 27776
rect 3315 27712 3331 27776
rect 3395 27712 3411 27776
rect 3475 27712 3483 27776
rect 3163 26688 3483 27712
rect 3163 26624 3171 26688
rect 3235 26624 3251 26688
rect 3315 26624 3331 26688
rect 3395 26624 3411 26688
rect 3475 26624 3483 26688
rect 3163 25600 3483 26624
rect 3163 25536 3171 25600
rect 3235 25536 3251 25600
rect 3315 25536 3331 25600
rect 3395 25536 3411 25600
rect 3475 25536 3483 25600
rect 3163 24512 3483 25536
rect 3163 24448 3171 24512
rect 3235 24448 3251 24512
rect 3315 24448 3331 24512
rect 3395 24448 3411 24512
rect 3475 24448 3483 24512
rect 3163 23424 3483 24448
rect 3163 23360 3171 23424
rect 3235 23360 3251 23424
rect 3315 23360 3331 23424
rect 3395 23360 3411 23424
rect 3475 23360 3483 23424
rect 3163 22336 3483 23360
rect 3163 22272 3171 22336
rect 3235 22272 3251 22336
rect 3315 22272 3331 22336
rect 3395 22272 3411 22336
rect 3475 22272 3483 22336
rect 3163 21248 3483 22272
rect 3163 21184 3171 21248
rect 3235 21184 3251 21248
rect 3315 21184 3331 21248
rect 3395 21184 3411 21248
rect 3475 21184 3483 21248
rect 3163 20160 3483 21184
rect 3163 20096 3171 20160
rect 3235 20096 3251 20160
rect 3315 20096 3331 20160
rect 3395 20096 3411 20160
rect 3475 20096 3483 20160
rect 3163 19072 3483 20096
rect 3163 19008 3171 19072
rect 3235 19008 3251 19072
rect 3315 19008 3331 19072
rect 3395 19008 3411 19072
rect 3475 19008 3483 19072
rect 3163 17984 3483 19008
rect 3163 17920 3171 17984
rect 3235 17920 3251 17984
rect 3315 17920 3331 17984
rect 3395 17920 3411 17984
rect 3475 17920 3483 17984
rect 3163 16896 3483 17920
rect 3163 16832 3171 16896
rect 3235 16832 3251 16896
rect 3315 16832 3331 16896
rect 3395 16832 3411 16896
rect 3475 16832 3483 16896
rect 3163 15808 3483 16832
rect 3163 15744 3171 15808
rect 3235 15744 3251 15808
rect 3315 15744 3331 15808
rect 3395 15744 3411 15808
rect 3475 15744 3483 15808
rect 3163 14720 3483 15744
rect 3163 14656 3171 14720
rect 3235 14656 3251 14720
rect 3315 14656 3331 14720
rect 3395 14656 3411 14720
rect 3475 14656 3483 14720
rect 3163 13632 3483 14656
rect 3163 13568 3171 13632
rect 3235 13568 3251 13632
rect 3315 13568 3331 13632
rect 3395 13568 3411 13632
rect 3475 13568 3483 13632
rect 3163 12544 3483 13568
rect 3163 12480 3171 12544
rect 3235 12480 3251 12544
rect 3315 12480 3331 12544
rect 3395 12480 3411 12544
rect 3475 12480 3483 12544
rect 3163 11456 3483 12480
rect 3163 11392 3171 11456
rect 3235 11392 3251 11456
rect 3315 11392 3331 11456
rect 3395 11392 3411 11456
rect 3475 11392 3483 11456
rect 3163 10368 3483 11392
rect 3163 10304 3171 10368
rect 3235 10304 3251 10368
rect 3315 10304 3331 10368
rect 3395 10304 3411 10368
rect 3475 10304 3483 10368
rect 3163 9280 3483 10304
rect 3163 9216 3171 9280
rect 3235 9216 3251 9280
rect 3315 9216 3331 9280
rect 3395 9216 3411 9280
rect 3475 9216 3483 9280
rect 3163 8192 3483 9216
rect 3163 8128 3171 8192
rect 3235 8128 3251 8192
rect 3315 8128 3331 8192
rect 3395 8128 3411 8192
rect 3475 8128 3483 8192
rect 3163 7104 3483 8128
rect 3163 7040 3171 7104
rect 3235 7040 3251 7104
rect 3315 7040 3331 7104
rect 3395 7040 3411 7104
rect 3475 7040 3483 7104
rect 3163 6016 3483 7040
rect 3163 5952 3171 6016
rect 3235 5952 3251 6016
rect 3315 5952 3331 6016
rect 3395 5952 3411 6016
rect 3475 5952 3483 6016
rect 3163 4928 3483 5952
rect 3163 4864 3171 4928
rect 3235 4864 3251 4928
rect 3315 4864 3331 4928
rect 3395 4864 3411 4928
rect 3475 4864 3483 4928
rect 3163 3840 3483 4864
rect 3163 3776 3171 3840
rect 3235 3776 3251 3840
rect 3315 3776 3331 3840
rect 3395 3776 3411 3840
rect 3475 3776 3483 3840
rect 3163 2752 3483 3776
rect 3163 2688 3171 2752
rect 3235 2688 3251 2752
rect 3315 2688 3331 2752
rect 3395 2688 3411 2752
rect 3475 2688 3483 2752
rect 3163 2128 3483 2688
rect 5382 46816 5702 47376
rect 5382 46752 5390 46816
rect 5454 46752 5470 46816
rect 5534 46752 5550 46816
rect 5614 46752 5630 46816
rect 5694 46752 5702 46816
rect 5382 45728 5702 46752
rect 5382 45664 5390 45728
rect 5454 45664 5470 45728
rect 5534 45664 5550 45728
rect 5614 45664 5630 45728
rect 5694 45664 5702 45728
rect 5382 44640 5702 45664
rect 5382 44576 5390 44640
rect 5454 44576 5470 44640
rect 5534 44576 5550 44640
rect 5614 44576 5630 44640
rect 5694 44576 5702 44640
rect 5382 43552 5702 44576
rect 5382 43488 5390 43552
rect 5454 43488 5470 43552
rect 5534 43488 5550 43552
rect 5614 43488 5630 43552
rect 5694 43488 5702 43552
rect 5382 42464 5702 43488
rect 5382 42400 5390 42464
rect 5454 42400 5470 42464
rect 5534 42400 5550 42464
rect 5614 42400 5630 42464
rect 5694 42400 5702 42464
rect 5382 41376 5702 42400
rect 5382 41312 5390 41376
rect 5454 41312 5470 41376
rect 5534 41312 5550 41376
rect 5614 41312 5630 41376
rect 5694 41312 5702 41376
rect 5382 40288 5702 41312
rect 5382 40224 5390 40288
rect 5454 40224 5470 40288
rect 5534 40224 5550 40288
rect 5614 40224 5630 40288
rect 5694 40224 5702 40288
rect 5382 39200 5702 40224
rect 5382 39136 5390 39200
rect 5454 39136 5470 39200
rect 5534 39136 5550 39200
rect 5614 39136 5630 39200
rect 5694 39136 5702 39200
rect 5382 38112 5702 39136
rect 5382 38048 5390 38112
rect 5454 38048 5470 38112
rect 5534 38048 5550 38112
rect 5614 38048 5630 38112
rect 5694 38048 5702 38112
rect 5382 37024 5702 38048
rect 5382 36960 5390 37024
rect 5454 36960 5470 37024
rect 5534 36960 5550 37024
rect 5614 36960 5630 37024
rect 5694 36960 5702 37024
rect 5382 35936 5702 36960
rect 5382 35872 5390 35936
rect 5454 35872 5470 35936
rect 5534 35872 5550 35936
rect 5614 35872 5630 35936
rect 5694 35872 5702 35936
rect 5382 34848 5702 35872
rect 5382 34784 5390 34848
rect 5454 34784 5470 34848
rect 5534 34784 5550 34848
rect 5614 34784 5630 34848
rect 5694 34784 5702 34848
rect 5382 33760 5702 34784
rect 5382 33696 5390 33760
rect 5454 33696 5470 33760
rect 5534 33696 5550 33760
rect 5614 33696 5630 33760
rect 5694 33696 5702 33760
rect 5382 32672 5702 33696
rect 5382 32608 5390 32672
rect 5454 32608 5470 32672
rect 5534 32608 5550 32672
rect 5614 32608 5630 32672
rect 5694 32608 5702 32672
rect 5382 31584 5702 32608
rect 5382 31520 5390 31584
rect 5454 31520 5470 31584
rect 5534 31520 5550 31584
rect 5614 31520 5630 31584
rect 5694 31520 5702 31584
rect 5382 30496 5702 31520
rect 5382 30432 5390 30496
rect 5454 30432 5470 30496
rect 5534 30432 5550 30496
rect 5614 30432 5630 30496
rect 5694 30432 5702 30496
rect 5382 29408 5702 30432
rect 5382 29344 5390 29408
rect 5454 29344 5470 29408
rect 5534 29344 5550 29408
rect 5614 29344 5630 29408
rect 5694 29344 5702 29408
rect 5382 28320 5702 29344
rect 5382 28256 5390 28320
rect 5454 28256 5470 28320
rect 5534 28256 5550 28320
rect 5614 28256 5630 28320
rect 5694 28256 5702 28320
rect 5382 27232 5702 28256
rect 5382 27168 5390 27232
rect 5454 27168 5470 27232
rect 5534 27168 5550 27232
rect 5614 27168 5630 27232
rect 5694 27168 5702 27232
rect 5382 26144 5702 27168
rect 5382 26080 5390 26144
rect 5454 26080 5470 26144
rect 5534 26080 5550 26144
rect 5614 26080 5630 26144
rect 5694 26080 5702 26144
rect 5382 25056 5702 26080
rect 5382 24992 5390 25056
rect 5454 24992 5470 25056
rect 5534 24992 5550 25056
rect 5614 24992 5630 25056
rect 5694 24992 5702 25056
rect 5382 23968 5702 24992
rect 5382 23904 5390 23968
rect 5454 23904 5470 23968
rect 5534 23904 5550 23968
rect 5614 23904 5630 23968
rect 5694 23904 5702 23968
rect 5382 22880 5702 23904
rect 5382 22816 5390 22880
rect 5454 22816 5470 22880
rect 5534 22816 5550 22880
rect 5614 22816 5630 22880
rect 5694 22816 5702 22880
rect 5382 21792 5702 22816
rect 5382 21728 5390 21792
rect 5454 21728 5470 21792
rect 5534 21728 5550 21792
rect 5614 21728 5630 21792
rect 5694 21728 5702 21792
rect 5382 20704 5702 21728
rect 5382 20640 5390 20704
rect 5454 20640 5470 20704
rect 5534 20640 5550 20704
rect 5614 20640 5630 20704
rect 5694 20640 5702 20704
rect 5382 19616 5702 20640
rect 5382 19552 5390 19616
rect 5454 19552 5470 19616
rect 5534 19552 5550 19616
rect 5614 19552 5630 19616
rect 5694 19552 5702 19616
rect 5382 18528 5702 19552
rect 5382 18464 5390 18528
rect 5454 18464 5470 18528
rect 5534 18464 5550 18528
rect 5614 18464 5630 18528
rect 5694 18464 5702 18528
rect 5382 17440 5702 18464
rect 5382 17376 5390 17440
rect 5454 17376 5470 17440
rect 5534 17376 5550 17440
rect 5614 17376 5630 17440
rect 5694 17376 5702 17440
rect 5382 16352 5702 17376
rect 5382 16288 5390 16352
rect 5454 16288 5470 16352
rect 5534 16288 5550 16352
rect 5614 16288 5630 16352
rect 5694 16288 5702 16352
rect 5382 15264 5702 16288
rect 5382 15200 5390 15264
rect 5454 15200 5470 15264
rect 5534 15200 5550 15264
rect 5614 15200 5630 15264
rect 5694 15200 5702 15264
rect 5382 14176 5702 15200
rect 5382 14112 5390 14176
rect 5454 14112 5470 14176
rect 5534 14112 5550 14176
rect 5614 14112 5630 14176
rect 5694 14112 5702 14176
rect 5382 13088 5702 14112
rect 5382 13024 5390 13088
rect 5454 13024 5470 13088
rect 5534 13024 5550 13088
rect 5614 13024 5630 13088
rect 5694 13024 5702 13088
rect 5382 12000 5702 13024
rect 5382 11936 5390 12000
rect 5454 11936 5470 12000
rect 5534 11936 5550 12000
rect 5614 11936 5630 12000
rect 5694 11936 5702 12000
rect 5382 10912 5702 11936
rect 5382 10848 5390 10912
rect 5454 10848 5470 10912
rect 5534 10848 5550 10912
rect 5614 10848 5630 10912
rect 5694 10848 5702 10912
rect 5382 9824 5702 10848
rect 5382 9760 5390 9824
rect 5454 9760 5470 9824
rect 5534 9760 5550 9824
rect 5614 9760 5630 9824
rect 5694 9760 5702 9824
rect 5382 8736 5702 9760
rect 5382 8672 5390 8736
rect 5454 8672 5470 8736
rect 5534 8672 5550 8736
rect 5614 8672 5630 8736
rect 5694 8672 5702 8736
rect 5382 7648 5702 8672
rect 5382 7584 5390 7648
rect 5454 7584 5470 7648
rect 5534 7584 5550 7648
rect 5614 7584 5630 7648
rect 5694 7584 5702 7648
rect 5382 6560 5702 7584
rect 5382 6496 5390 6560
rect 5454 6496 5470 6560
rect 5534 6496 5550 6560
rect 5614 6496 5630 6560
rect 5694 6496 5702 6560
rect 5382 5472 5702 6496
rect 5382 5408 5390 5472
rect 5454 5408 5470 5472
rect 5534 5408 5550 5472
rect 5614 5408 5630 5472
rect 5694 5408 5702 5472
rect 5382 4384 5702 5408
rect 5382 4320 5390 4384
rect 5454 4320 5470 4384
rect 5534 4320 5550 4384
rect 5614 4320 5630 4384
rect 5694 4320 5702 4384
rect 5382 3296 5702 4320
rect 5382 3232 5390 3296
rect 5454 3232 5470 3296
rect 5534 3232 5550 3296
rect 5614 3232 5630 3296
rect 5694 3232 5702 3296
rect 5382 2208 5702 3232
rect 5382 2144 5390 2208
rect 5454 2144 5470 2208
rect 5534 2144 5550 2208
rect 5614 2144 5630 2208
rect 5694 2144 5702 2208
rect 5382 2128 5702 2144
rect 7602 47360 7922 47376
rect 7602 47296 7610 47360
rect 7674 47296 7690 47360
rect 7754 47296 7770 47360
rect 7834 47296 7850 47360
rect 7914 47296 7922 47360
rect 7602 46272 7922 47296
rect 7602 46208 7610 46272
rect 7674 46208 7690 46272
rect 7754 46208 7770 46272
rect 7834 46208 7850 46272
rect 7914 46208 7922 46272
rect 7602 45184 7922 46208
rect 7602 45120 7610 45184
rect 7674 45120 7690 45184
rect 7754 45120 7770 45184
rect 7834 45120 7850 45184
rect 7914 45120 7922 45184
rect 7602 44096 7922 45120
rect 7602 44032 7610 44096
rect 7674 44032 7690 44096
rect 7754 44032 7770 44096
rect 7834 44032 7850 44096
rect 7914 44032 7922 44096
rect 7602 43008 7922 44032
rect 7602 42944 7610 43008
rect 7674 42944 7690 43008
rect 7754 42944 7770 43008
rect 7834 42944 7850 43008
rect 7914 42944 7922 43008
rect 7602 41920 7922 42944
rect 7602 41856 7610 41920
rect 7674 41856 7690 41920
rect 7754 41856 7770 41920
rect 7834 41856 7850 41920
rect 7914 41856 7922 41920
rect 7602 40832 7922 41856
rect 7602 40768 7610 40832
rect 7674 40768 7690 40832
rect 7754 40768 7770 40832
rect 7834 40768 7850 40832
rect 7914 40768 7922 40832
rect 7602 39744 7922 40768
rect 7602 39680 7610 39744
rect 7674 39680 7690 39744
rect 7754 39680 7770 39744
rect 7834 39680 7850 39744
rect 7914 39680 7922 39744
rect 7602 38656 7922 39680
rect 7602 38592 7610 38656
rect 7674 38592 7690 38656
rect 7754 38592 7770 38656
rect 7834 38592 7850 38656
rect 7914 38592 7922 38656
rect 7602 37568 7922 38592
rect 7602 37504 7610 37568
rect 7674 37504 7690 37568
rect 7754 37504 7770 37568
rect 7834 37504 7850 37568
rect 7914 37504 7922 37568
rect 7602 36480 7922 37504
rect 7602 36416 7610 36480
rect 7674 36416 7690 36480
rect 7754 36416 7770 36480
rect 7834 36416 7850 36480
rect 7914 36416 7922 36480
rect 7602 35392 7922 36416
rect 7602 35328 7610 35392
rect 7674 35328 7690 35392
rect 7754 35328 7770 35392
rect 7834 35328 7850 35392
rect 7914 35328 7922 35392
rect 7602 34304 7922 35328
rect 7602 34240 7610 34304
rect 7674 34240 7690 34304
rect 7754 34240 7770 34304
rect 7834 34240 7850 34304
rect 7914 34240 7922 34304
rect 7602 33216 7922 34240
rect 7602 33152 7610 33216
rect 7674 33152 7690 33216
rect 7754 33152 7770 33216
rect 7834 33152 7850 33216
rect 7914 33152 7922 33216
rect 7602 32128 7922 33152
rect 7602 32064 7610 32128
rect 7674 32064 7690 32128
rect 7754 32064 7770 32128
rect 7834 32064 7850 32128
rect 7914 32064 7922 32128
rect 7602 31040 7922 32064
rect 7602 30976 7610 31040
rect 7674 30976 7690 31040
rect 7754 30976 7770 31040
rect 7834 30976 7850 31040
rect 7914 30976 7922 31040
rect 7602 29952 7922 30976
rect 7602 29888 7610 29952
rect 7674 29888 7690 29952
rect 7754 29888 7770 29952
rect 7834 29888 7850 29952
rect 7914 29888 7922 29952
rect 7602 28864 7922 29888
rect 7602 28800 7610 28864
rect 7674 28800 7690 28864
rect 7754 28800 7770 28864
rect 7834 28800 7850 28864
rect 7914 28800 7922 28864
rect 7602 27776 7922 28800
rect 7602 27712 7610 27776
rect 7674 27712 7690 27776
rect 7754 27712 7770 27776
rect 7834 27712 7850 27776
rect 7914 27712 7922 27776
rect 7602 26688 7922 27712
rect 7602 26624 7610 26688
rect 7674 26624 7690 26688
rect 7754 26624 7770 26688
rect 7834 26624 7850 26688
rect 7914 26624 7922 26688
rect 7602 25600 7922 26624
rect 7602 25536 7610 25600
rect 7674 25536 7690 25600
rect 7754 25536 7770 25600
rect 7834 25536 7850 25600
rect 7914 25536 7922 25600
rect 7602 24512 7922 25536
rect 7602 24448 7610 24512
rect 7674 24448 7690 24512
rect 7754 24448 7770 24512
rect 7834 24448 7850 24512
rect 7914 24448 7922 24512
rect 7602 23424 7922 24448
rect 7602 23360 7610 23424
rect 7674 23360 7690 23424
rect 7754 23360 7770 23424
rect 7834 23360 7850 23424
rect 7914 23360 7922 23424
rect 7602 22336 7922 23360
rect 7602 22272 7610 22336
rect 7674 22272 7690 22336
rect 7754 22272 7770 22336
rect 7834 22272 7850 22336
rect 7914 22272 7922 22336
rect 7602 21248 7922 22272
rect 7602 21184 7610 21248
rect 7674 21184 7690 21248
rect 7754 21184 7770 21248
rect 7834 21184 7850 21248
rect 7914 21184 7922 21248
rect 7602 20160 7922 21184
rect 7602 20096 7610 20160
rect 7674 20096 7690 20160
rect 7754 20096 7770 20160
rect 7834 20096 7850 20160
rect 7914 20096 7922 20160
rect 7602 19072 7922 20096
rect 7602 19008 7610 19072
rect 7674 19008 7690 19072
rect 7754 19008 7770 19072
rect 7834 19008 7850 19072
rect 7914 19008 7922 19072
rect 7602 17984 7922 19008
rect 7602 17920 7610 17984
rect 7674 17920 7690 17984
rect 7754 17920 7770 17984
rect 7834 17920 7850 17984
rect 7914 17920 7922 17984
rect 7602 16896 7922 17920
rect 7602 16832 7610 16896
rect 7674 16832 7690 16896
rect 7754 16832 7770 16896
rect 7834 16832 7850 16896
rect 7914 16832 7922 16896
rect 7602 15808 7922 16832
rect 7602 15744 7610 15808
rect 7674 15744 7690 15808
rect 7754 15744 7770 15808
rect 7834 15744 7850 15808
rect 7914 15744 7922 15808
rect 7602 14720 7922 15744
rect 7602 14656 7610 14720
rect 7674 14656 7690 14720
rect 7754 14656 7770 14720
rect 7834 14656 7850 14720
rect 7914 14656 7922 14720
rect 7602 13632 7922 14656
rect 7602 13568 7610 13632
rect 7674 13568 7690 13632
rect 7754 13568 7770 13632
rect 7834 13568 7850 13632
rect 7914 13568 7922 13632
rect 7602 12544 7922 13568
rect 7602 12480 7610 12544
rect 7674 12480 7690 12544
rect 7754 12480 7770 12544
rect 7834 12480 7850 12544
rect 7914 12480 7922 12544
rect 7602 11456 7922 12480
rect 7602 11392 7610 11456
rect 7674 11392 7690 11456
rect 7754 11392 7770 11456
rect 7834 11392 7850 11456
rect 7914 11392 7922 11456
rect 7602 10368 7922 11392
rect 7602 10304 7610 10368
rect 7674 10304 7690 10368
rect 7754 10304 7770 10368
rect 7834 10304 7850 10368
rect 7914 10304 7922 10368
rect 7602 9280 7922 10304
rect 7602 9216 7610 9280
rect 7674 9216 7690 9280
rect 7754 9216 7770 9280
rect 7834 9216 7850 9280
rect 7914 9216 7922 9280
rect 7602 8192 7922 9216
rect 7602 8128 7610 8192
rect 7674 8128 7690 8192
rect 7754 8128 7770 8192
rect 7834 8128 7850 8192
rect 7914 8128 7922 8192
rect 7602 7104 7922 8128
rect 7602 7040 7610 7104
rect 7674 7040 7690 7104
rect 7754 7040 7770 7104
rect 7834 7040 7850 7104
rect 7914 7040 7922 7104
rect 7602 6016 7922 7040
rect 7602 5952 7610 6016
rect 7674 5952 7690 6016
rect 7754 5952 7770 6016
rect 7834 5952 7850 6016
rect 7914 5952 7922 6016
rect 7602 4928 7922 5952
rect 7602 4864 7610 4928
rect 7674 4864 7690 4928
rect 7754 4864 7770 4928
rect 7834 4864 7850 4928
rect 7914 4864 7922 4928
rect 7602 3840 7922 4864
rect 7602 3776 7610 3840
rect 7674 3776 7690 3840
rect 7754 3776 7770 3840
rect 7834 3776 7850 3840
rect 7914 3776 7922 3840
rect 7602 2752 7922 3776
rect 7602 2688 7610 2752
rect 7674 2688 7690 2752
rect 7754 2688 7770 2752
rect 7834 2688 7850 2752
rect 7914 2688 7922 2752
rect 7602 2128 7922 2688
rect 9821 46816 10141 47376
rect 9821 46752 9829 46816
rect 9893 46752 9909 46816
rect 9973 46752 9989 46816
rect 10053 46752 10069 46816
rect 10133 46752 10141 46816
rect 9821 45728 10141 46752
rect 9821 45664 9829 45728
rect 9893 45664 9909 45728
rect 9973 45664 9989 45728
rect 10053 45664 10069 45728
rect 10133 45664 10141 45728
rect 9821 44640 10141 45664
rect 9821 44576 9829 44640
rect 9893 44576 9909 44640
rect 9973 44576 9989 44640
rect 10053 44576 10069 44640
rect 10133 44576 10141 44640
rect 9821 43552 10141 44576
rect 9821 43488 9829 43552
rect 9893 43488 9909 43552
rect 9973 43488 9989 43552
rect 10053 43488 10069 43552
rect 10133 43488 10141 43552
rect 9821 42464 10141 43488
rect 9821 42400 9829 42464
rect 9893 42400 9909 42464
rect 9973 42400 9989 42464
rect 10053 42400 10069 42464
rect 10133 42400 10141 42464
rect 9821 41376 10141 42400
rect 9821 41312 9829 41376
rect 9893 41312 9909 41376
rect 9973 41312 9989 41376
rect 10053 41312 10069 41376
rect 10133 41312 10141 41376
rect 9821 40288 10141 41312
rect 9821 40224 9829 40288
rect 9893 40224 9909 40288
rect 9973 40224 9989 40288
rect 10053 40224 10069 40288
rect 10133 40224 10141 40288
rect 9821 39200 10141 40224
rect 9821 39136 9829 39200
rect 9893 39136 9909 39200
rect 9973 39136 9989 39200
rect 10053 39136 10069 39200
rect 10133 39136 10141 39200
rect 9821 38112 10141 39136
rect 9821 38048 9829 38112
rect 9893 38048 9909 38112
rect 9973 38048 9989 38112
rect 10053 38048 10069 38112
rect 10133 38048 10141 38112
rect 9821 37024 10141 38048
rect 9821 36960 9829 37024
rect 9893 36960 9909 37024
rect 9973 36960 9989 37024
rect 10053 36960 10069 37024
rect 10133 36960 10141 37024
rect 9821 35936 10141 36960
rect 9821 35872 9829 35936
rect 9893 35872 9909 35936
rect 9973 35872 9989 35936
rect 10053 35872 10069 35936
rect 10133 35872 10141 35936
rect 9821 34848 10141 35872
rect 9821 34784 9829 34848
rect 9893 34784 9909 34848
rect 9973 34784 9989 34848
rect 10053 34784 10069 34848
rect 10133 34784 10141 34848
rect 9821 33760 10141 34784
rect 9821 33696 9829 33760
rect 9893 33696 9909 33760
rect 9973 33696 9989 33760
rect 10053 33696 10069 33760
rect 10133 33696 10141 33760
rect 9821 32672 10141 33696
rect 9821 32608 9829 32672
rect 9893 32608 9909 32672
rect 9973 32608 9989 32672
rect 10053 32608 10069 32672
rect 10133 32608 10141 32672
rect 9821 31584 10141 32608
rect 9821 31520 9829 31584
rect 9893 31520 9909 31584
rect 9973 31520 9989 31584
rect 10053 31520 10069 31584
rect 10133 31520 10141 31584
rect 9821 30496 10141 31520
rect 9821 30432 9829 30496
rect 9893 30432 9909 30496
rect 9973 30432 9989 30496
rect 10053 30432 10069 30496
rect 10133 30432 10141 30496
rect 9821 29408 10141 30432
rect 9821 29344 9829 29408
rect 9893 29344 9909 29408
rect 9973 29344 9989 29408
rect 10053 29344 10069 29408
rect 10133 29344 10141 29408
rect 9821 28320 10141 29344
rect 9821 28256 9829 28320
rect 9893 28256 9909 28320
rect 9973 28256 9989 28320
rect 10053 28256 10069 28320
rect 10133 28256 10141 28320
rect 9821 27232 10141 28256
rect 9821 27168 9829 27232
rect 9893 27168 9909 27232
rect 9973 27168 9989 27232
rect 10053 27168 10069 27232
rect 10133 27168 10141 27232
rect 9821 26144 10141 27168
rect 9821 26080 9829 26144
rect 9893 26080 9909 26144
rect 9973 26080 9989 26144
rect 10053 26080 10069 26144
rect 10133 26080 10141 26144
rect 9821 25056 10141 26080
rect 9821 24992 9829 25056
rect 9893 24992 9909 25056
rect 9973 24992 9989 25056
rect 10053 24992 10069 25056
rect 10133 24992 10141 25056
rect 9821 23968 10141 24992
rect 9821 23904 9829 23968
rect 9893 23904 9909 23968
rect 9973 23904 9989 23968
rect 10053 23904 10069 23968
rect 10133 23904 10141 23968
rect 9821 22880 10141 23904
rect 9821 22816 9829 22880
rect 9893 22816 9909 22880
rect 9973 22816 9989 22880
rect 10053 22816 10069 22880
rect 10133 22816 10141 22880
rect 9821 21792 10141 22816
rect 9821 21728 9829 21792
rect 9893 21728 9909 21792
rect 9973 21728 9989 21792
rect 10053 21728 10069 21792
rect 10133 21728 10141 21792
rect 9821 20704 10141 21728
rect 9821 20640 9829 20704
rect 9893 20640 9909 20704
rect 9973 20640 9989 20704
rect 10053 20640 10069 20704
rect 10133 20640 10141 20704
rect 9821 19616 10141 20640
rect 9821 19552 9829 19616
rect 9893 19552 9909 19616
rect 9973 19552 9989 19616
rect 10053 19552 10069 19616
rect 10133 19552 10141 19616
rect 9821 18528 10141 19552
rect 9821 18464 9829 18528
rect 9893 18464 9909 18528
rect 9973 18464 9989 18528
rect 10053 18464 10069 18528
rect 10133 18464 10141 18528
rect 9821 17440 10141 18464
rect 9821 17376 9829 17440
rect 9893 17376 9909 17440
rect 9973 17376 9989 17440
rect 10053 17376 10069 17440
rect 10133 17376 10141 17440
rect 9821 16352 10141 17376
rect 9821 16288 9829 16352
rect 9893 16288 9909 16352
rect 9973 16288 9989 16352
rect 10053 16288 10069 16352
rect 10133 16288 10141 16352
rect 9821 15264 10141 16288
rect 9821 15200 9829 15264
rect 9893 15200 9909 15264
rect 9973 15200 9989 15264
rect 10053 15200 10069 15264
rect 10133 15200 10141 15264
rect 9821 14176 10141 15200
rect 9821 14112 9829 14176
rect 9893 14112 9909 14176
rect 9973 14112 9989 14176
rect 10053 14112 10069 14176
rect 10133 14112 10141 14176
rect 9821 13088 10141 14112
rect 9821 13024 9829 13088
rect 9893 13024 9909 13088
rect 9973 13024 9989 13088
rect 10053 13024 10069 13088
rect 10133 13024 10141 13088
rect 9821 12000 10141 13024
rect 9821 11936 9829 12000
rect 9893 11936 9909 12000
rect 9973 11936 9989 12000
rect 10053 11936 10069 12000
rect 10133 11936 10141 12000
rect 9821 10912 10141 11936
rect 9821 10848 9829 10912
rect 9893 10848 9909 10912
rect 9973 10848 9989 10912
rect 10053 10848 10069 10912
rect 10133 10848 10141 10912
rect 9821 9824 10141 10848
rect 9821 9760 9829 9824
rect 9893 9760 9909 9824
rect 9973 9760 9989 9824
rect 10053 9760 10069 9824
rect 10133 9760 10141 9824
rect 9821 8736 10141 9760
rect 9821 8672 9829 8736
rect 9893 8672 9909 8736
rect 9973 8672 9989 8736
rect 10053 8672 10069 8736
rect 10133 8672 10141 8736
rect 9821 7648 10141 8672
rect 9821 7584 9829 7648
rect 9893 7584 9909 7648
rect 9973 7584 9989 7648
rect 10053 7584 10069 7648
rect 10133 7584 10141 7648
rect 9821 6560 10141 7584
rect 9821 6496 9829 6560
rect 9893 6496 9909 6560
rect 9973 6496 9989 6560
rect 10053 6496 10069 6560
rect 10133 6496 10141 6560
rect 9821 5472 10141 6496
rect 9821 5408 9829 5472
rect 9893 5408 9909 5472
rect 9973 5408 9989 5472
rect 10053 5408 10069 5472
rect 10133 5408 10141 5472
rect 9821 4384 10141 5408
rect 9821 4320 9829 4384
rect 9893 4320 9909 4384
rect 9973 4320 9989 4384
rect 10053 4320 10069 4384
rect 10133 4320 10141 4384
rect 9821 3296 10141 4320
rect 9821 3232 9829 3296
rect 9893 3232 9909 3296
rect 9973 3232 9989 3296
rect 10053 3232 10069 3296
rect 10133 3232 10141 3296
rect 9821 2208 10141 3232
rect 9821 2144 9829 2208
rect 9893 2144 9909 2208
rect 9973 2144 9989 2208
rect 10053 2144 10069 2208
rect 10133 2144 10141 2208
rect 9821 2128 10141 2144
rect 12041 47360 12361 47376
rect 12041 47296 12049 47360
rect 12113 47296 12129 47360
rect 12193 47296 12209 47360
rect 12273 47296 12289 47360
rect 12353 47296 12361 47360
rect 12041 46272 12361 47296
rect 12041 46208 12049 46272
rect 12113 46208 12129 46272
rect 12193 46208 12209 46272
rect 12273 46208 12289 46272
rect 12353 46208 12361 46272
rect 12041 45184 12361 46208
rect 12041 45120 12049 45184
rect 12113 45120 12129 45184
rect 12193 45120 12209 45184
rect 12273 45120 12289 45184
rect 12353 45120 12361 45184
rect 12041 44096 12361 45120
rect 12041 44032 12049 44096
rect 12113 44032 12129 44096
rect 12193 44032 12209 44096
rect 12273 44032 12289 44096
rect 12353 44032 12361 44096
rect 12041 43008 12361 44032
rect 12041 42944 12049 43008
rect 12113 42944 12129 43008
rect 12193 42944 12209 43008
rect 12273 42944 12289 43008
rect 12353 42944 12361 43008
rect 12041 41920 12361 42944
rect 12041 41856 12049 41920
rect 12113 41856 12129 41920
rect 12193 41856 12209 41920
rect 12273 41856 12289 41920
rect 12353 41856 12361 41920
rect 12041 40832 12361 41856
rect 12041 40768 12049 40832
rect 12113 40768 12129 40832
rect 12193 40768 12209 40832
rect 12273 40768 12289 40832
rect 12353 40768 12361 40832
rect 12041 39744 12361 40768
rect 12041 39680 12049 39744
rect 12113 39680 12129 39744
rect 12193 39680 12209 39744
rect 12273 39680 12289 39744
rect 12353 39680 12361 39744
rect 12041 38656 12361 39680
rect 12041 38592 12049 38656
rect 12113 38592 12129 38656
rect 12193 38592 12209 38656
rect 12273 38592 12289 38656
rect 12353 38592 12361 38656
rect 12041 37568 12361 38592
rect 12041 37504 12049 37568
rect 12113 37504 12129 37568
rect 12193 37504 12209 37568
rect 12273 37504 12289 37568
rect 12353 37504 12361 37568
rect 12041 36480 12361 37504
rect 12041 36416 12049 36480
rect 12113 36416 12129 36480
rect 12193 36416 12209 36480
rect 12273 36416 12289 36480
rect 12353 36416 12361 36480
rect 12041 35392 12361 36416
rect 12041 35328 12049 35392
rect 12113 35328 12129 35392
rect 12193 35328 12209 35392
rect 12273 35328 12289 35392
rect 12353 35328 12361 35392
rect 12041 34304 12361 35328
rect 12041 34240 12049 34304
rect 12113 34240 12129 34304
rect 12193 34240 12209 34304
rect 12273 34240 12289 34304
rect 12353 34240 12361 34304
rect 12041 33216 12361 34240
rect 12041 33152 12049 33216
rect 12113 33152 12129 33216
rect 12193 33152 12209 33216
rect 12273 33152 12289 33216
rect 12353 33152 12361 33216
rect 12041 32128 12361 33152
rect 12041 32064 12049 32128
rect 12113 32064 12129 32128
rect 12193 32064 12209 32128
rect 12273 32064 12289 32128
rect 12353 32064 12361 32128
rect 12041 31040 12361 32064
rect 12041 30976 12049 31040
rect 12113 30976 12129 31040
rect 12193 30976 12209 31040
rect 12273 30976 12289 31040
rect 12353 30976 12361 31040
rect 12041 29952 12361 30976
rect 12041 29888 12049 29952
rect 12113 29888 12129 29952
rect 12193 29888 12209 29952
rect 12273 29888 12289 29952
rect 12353 29888 12361 29952
rect 12041 28864 12361 29888
rect 12041 28800 12049 28864
rect 12113 28800 12129 28864
rect 12193 28800 12209 28864
rect 12273 28800 12289 28864
rect 12353 28800 12361 28864
rect 12041 27776 12361 28800
rect 12041 27712 12049 27776
rect 12113 27712 12129 27776
rect 12193 27712 12209 27776
rect 12273 27712 12289 27776
rect 12353 27712 12361 27776
rect 12041 26688 12361 27712
rect 12041 26624 12049 26688
rect 12113 26624 12129 26688
rect 12193 26624 12209 26688
rect 12273 26624 12289 26688
rect 12353 26624 12361 26688
rect 12041 25600 12361 26624
rect 12041 25536 12049 25600
rect 12113 25536 12129 25600
rect 12193 25536 12209 25600
rect 12273 25536 12289 25600
rect 12353 25536 12361 25600
rect 12041 24512 12361 25536
rect 12041 24448 12049 24512
rect 12113 24448 12129 24512
rect 12193 24448 12209 24512
rect 12273 24448 12289 24512
rect 12353 24448 12361 24512
rect 12041 23424 12361 24448
rect 12041 23360 12049 23424
rect 12113 23360 12129 23424
rect 12193 23360 12209 23424
rect 12273 23360 12289 23424
rect 12353 23360 12361 23424
rect 12041 22336 12361 23360
rect 12041 22272 12049 22336
rect 12113 22272 12129 22336
rect 12193 22272 12209 22336
rect 12273 22272 12289 22336
rect 12353 22272 12361 22336
rect 12041 21248 12361 22272
rect 12041 21184 12049 21248
rect 12113 21184 12129 21248
rect 12193 21184 12209 21248
rect 12273 21184 12289 21248
rect 12353 21184 12361 21248
rect 12041 20160 12361 21184
rect 12041 20096 12049 20160
rect 12113 20096 12129 20160
rect 12193 20096 12209 20160
rect 12273 20096 12289 20160
rect 12353 20096 12361 20160
rect 12041 19072 12361 20096
rect 12041 19008 12049 19072
rect 12113 19008 12129 19072
rect 12193 19008 12209 19072
rect 12273 19008 12289 19072
rect 12353 19008 12361 19072
rect 12041 17984 12361 19008
rect 12041 17920 12049 17984
rect 12113 17920 12129 17984
rect 12193 17920 12209 17984
rect 12273 17920 12289 17984
rect 12353 17920 12361 17984
rect 12041 16896 12361 17920
rect 12041 16832 12049 16896
rect 12113 16832 12129 16896
rect 12193 16832 12209 16896
rect 12273 16832 12289 16896
rect 12353 16832 12361 16896
rect 12041 15808 12361 16832
rect 12041 15744 12049 15808
rect 12113 15744 12129 15808
rect 12193 15744 12209 15808
rect 12273 15744 12289 15808
rect 12353 15744 12361 15808
rect 12041 14720 12361 15744
rect 12041 14656 12049 14720
rect 12113 14656 12129 14720
rect 12193 14656 12209 14720
rect 12273 14656 12289 14720
rect 12353 14656 12361 14720
rect 12041 13632 12361 14656
rect 12041 13568 12049 13632
rect 12113 13568 12129 13632
rect 12193 13568 12209 13632
rect 12273 13568 12289 13632
rect 12353 13568 12361 13632
rect 12041 12544 12361 13568
rect 12041 12480 12049 12544
rect 12113 12480 12129 12544
rect 12193 12480 12209 12544
rect 12273 12480 12289 12544
rect 12353 12480 12361 12544
rect 12041 11456 12361 12480
rect 12041 11392 12049 11456
rect 12113 11392 12129 11456
rect 12193 11392 12209 11456
rect 12273 11392 12289 11456
rect 12353 11392 12361 11456
rect 12041 10368 12361 11392
rect 12041 10304 12049 10368
rect 12113 10304 12129 10368
rect 12193 10304 12209 10368
rect 12273 10304 12289 10368
rect 12353 10304 12361 10368
rect 12041 9280 12361 10304
rect 12041 9216 12049 9280
rect 12113 9216 12129 9280
rect 12193 9216 12209 9280
rect 12273 9216 12289 9280
rect 12353 9216 12361 9280
rect 12041 8192 12361 9216
rect 12041 8128 12049 8192
rect 12113 8128 12129 8192
rect 12193 8128 12209 8192
rect 12273 8128 12289 8192
rect 12353 8128 12361 8192
rect 12041 7104 12361 8128
rect 12041 7040 12049 7104
rect 12113 7040 12129 7104
rect 12193 7040 12209 7104
rect 12273 7040 12289 7104
rect 12353 7040 12361 7104
rect 12041 6016 12361 7040
rect 12041 5952 12049 6016
rect 12113 5952 12129 6016
rect 12193 5952 12209 6016
rect 12273 5952 12289 6016
rect 12353 5952 12361 6016
rect 12041 4928 12361 5952
rect 12041 4864 12049 4928
rect 12113 4864 12129 4928
rect 12193 4864 12209 4928
rect 12273 4864 12289 4928
rect 12353 4864 12361 4928
rect 12041 3840 12361 4864
rect 12041 3776 12049 3840
rect 12113 3776 12129 3840
rect 12193 3776 12209 3840
rect 12273 3776 12289 3840
rect 12353 3776 12361 3840
rect 12041 2752 12361 3776
rect 12041 2688 12049 2752
rect 12113 2688 12129 2752
rect 12193 2688 12209 2752
rect 12273 2688 12289 2752
rect 12353 2688 12361 2752
rect 12041 2128 12361 2688
rect 14260 46816 14580 47376
rect 14260 46752 14268 46816
rect 14332 46752 14348 46816
rect 14412 46752 14428 46816
rect 14492 46752 14508 46816
rect 14572 46752 14580 46816
rect 14260 45728 14580 46752
rect 14260 45664 14268 45728
rect 14332 45664 14348 45728
rect 14412 45664 14428 45728
rect 14492 45664 14508 45728
rect 14572 45664 14580 45728
rect 14260 44640 14580 45664
rect 14260 44576 14268 44640
rect 14332 44576 14348 44640
rect 14412 44576 14428 44640
rect 14492 44576 14508 44640
rect 14572 44576 14580 44640
rect 14260 43552 14580 44576
rect 14260 43488 14268 43552
rect 14332 43488 14348 43552
rect 14412 43488 14428 43552
rect 14492 43488 14508 43552
rect 14572 43488 14580 43552
rect 14260 42464 14580 43488
rect 14260 42400 14268 42464
rect 14332 42400 14348 42464
rect 14412 42400 14428 42464
rect 14492 42400 14508 42464
rect 14572 42400 14580 42464
rect 14260 41376 14580 42400
rect 14260 41312 14268 41376
rect 14332 41312 14348 41376
rect 14412 41312 14428 41376
rect 14492 41312 14508 41376
rect 14572 41312 14580 41376
rect 14260 40288 14580 41312
rect 14260 40224 14268 40288
rect 14332 40224 14348 40288
rect 14412 40224 14428 40288
rect 14492 40224 14508 40288
rect 14572 40224 14580 40288
rect 14260 39200 14580 40224
rect 14260 39136 14268 39200
rect 14332 39136 14348 39200
rect 14412 39136 14428 39200
rect 14492 39136 14508 39200
rect 14572 39136 14580 39200
rect 14260 38112 14580 39136
rect 14260 38048 14268 38112
rect 14332 38048 14348 38112
rect 14412 38048 14428 38112
rect 14492 38048 14508 38112
rect 14572 38048 14580 38112
rect 14260 37024 14580 38048
rect 14260 36960 14268 37024
rect 14332 36960 14348 37024
rect 14412 36960 14428 37024
rect 14492 36960 14508 37024
rect 14572 36960 14580 37024
rect 14260 35936 14580 36960
rect 14260 35872 14268 35936
rect 14332 35872 14348 35936
rect 14412 35872 14428 35936
rect 14492 35872 14508 35936
rect 14572 35872 14580 35936
rect 14260 34848 14580 35872
rect 14260 34784 14268 34848
rect 14332 34784 14348 34848
rect 14412 34784 14428 34848
rect 14492 34784 14508 34848
rect 14572 34784 14580 34848
rect 14260 33760 14580 34784
rect 14260 33696 14268 33760
rect 14332 33696 14348 33760
rect 14412 33696 14428 33760
rect 14492 33696 14508 33760
rect 14572 33696 14580 33760
rect 14260 32672 14580 33696
rect 14260 32608 14268 32672
rect 14332 32608 14348 32672
rect 14412 32608 14428 32672
rect 14492 32608 14508 32672
rect 14572 32608 14580 32672
rect 14260 31584 14580 32608
rect 14260 31520 14268 31584
rect 14332 31520 14348 31584
rect 14412 31520 14428 31584
rect 14492 31520 14508 31584
rect 14572 31520 14580 31584
rect 14260 30496 14580 31520
rect 14260 30432 14268 30496
rect 14332 30432 14348 30496
rect 14412 30432 14428 30496
rect 14492 30432 14508 30496
rect 14572 30432 14580 30496
rect 14260 29408 14580 30432
rect 14260 29344 14268 29408
rect 14332 29344 14348 29408
rect 14412 29344 14428 29408
rect 14492 29344 14508 29408
rect 14572 29344 14580 29408
rect 14260 28320 14580 29344
rect 14260 28256 14268 28320
rect 14332 28256 14348 28320
rect 14412 28256 14428 28320
rect 14492 28256 14508 28320
rect 14572 28256 14580 28320
rect 14260 27232 14580 28256
rect 14260 27168 14268 27232
rect 14332 27168 14348 27232
rect 14412 27168 14428 27232
rect 14492 27168 14508 27232
rect 14572 27168 14580 27232
rect 14260 26144 14580 27168
rect 14260 26080 14268 26144
rect 14332 26080 14348 26144
rect 14412 26080 14428 26144
rect 14492 26080 14508 26144
rect 14572 26080 14580 26144
rect 14260 25056 14580 26080
rect 14260 24992 14268 25056
rect 14332 24992 14348 25056
rect 14412 24992 14428 25056
rect 14492 24992 14508 25056
rect 14572 24992 14580 25056
rect 14260 23968 14580 24992
rect 14260 23904 14268 23968
rect 14332 23904 14348 23968
rect 14412 23904 14428 23968
rect 14492 23904 14508 23968
rect 14572 23904 14580 23968
rect 14260 22880 14580 23904
rect 14260 22816 14268 22880
rect 14332 22816 14348 22880
rect 14412 22816 14428 22880
rect 14492 22816 14508 22880
rect 14572 22816 14580 22880
rect 14260 21792 14580 22816
rect 14260 21728 14268 21792
rect 14332 21728 14348 21792
rect 14412 21728 14428 21792
rect 14492 21728 14508 21792
rect 14572 21728 14580 21792
rect 14260 20704 14580 21728
rect 14260 20640 14268 20704
rect 14332 20640 14348 20704
rect 14412 20640 14428 20704
rect 14492 20640 14508 20704
rect 14572 20640 14580 20704
rect 14260 19616 14580 20640
rect 14260 19552 14268 19616
rect 14332 19552 14348 19616
rect 14412 19552 14428 19616
rect 14492 19552 14508 19616
rect 14572 19552 14580 19616
rect 14260 18528 14580 19552
rect 14260 18464 14268 18528
rect 14332 18464 14348 18528
rect 14412 18464 14428 18528
rect 14492 18464 14508 18528
rect 14572 18464 14580 18528
rect 14260 17440 14580 18464
rect 14260 17376 14268 17440
rect 14332 17376 14348 17440
rect 14412 17376 14428 17440
rect 14492 17376 14508 17440
rect 14572 17376 14580 17440
rect 14260 16352 14580 17376
rect 14260 16288 14268 16352
rect 14332 16288 14348 16352
rect 14412 16288 14428 16352
rect 14492 16288 14508 16352
rect 14572 16288 14580 16352
rect 14260 15264 14580 16288
rect 14260 15200 14268 15264
rect 14332 15200 14348 15264
rect 14412 15200 14428 15264
rect 14492 15200 14508 15264
rect 14572 15200 14580 15264
rect 14260 14176 14580 15200
rect 14260 14112 14268 14176
rect 14332 14112 14348 14176
rect 14412 14112 14428 14176
rect 14492 14112 14508 14176
rect 14572 14112 14580 14176
rect 14260 13088 14580 14112
rect 14260 13024 14268 13088
rect 14332 13024 14348 13088
rect 14412 13024 14428 13088
rect 14492 13024 14508 13088
rect 14572 13024 14580 13088
rect 14260 12000 14580 13024
rect 14260 11936 14268 12000
rect 14332 11936 14348 12000
rect 14412 11936 14428 12000
rect 14492 11936 14508 12000
rect 14572 11936 14580 12000
rect 14260 10912 14580 11936
rect 14260 10848 14268 10912
rect 14332 10848 14348 10912
rect 14412 10848 14428 10912
rect 14492 10848 14508 10912
rect 14572 10848 14580 10912
rect 14260 9824 14580 10848
rect 14260 9760 14268 9824
rect 14332 9760 14348 9824
rect 14412 9760 14428 9824
rect 14492 9760 14508 9824
rect 14572 9760 14580 9824
rect 14260 8736 14580 9760
rect 14260 8672 14268 8736
rect 14332 8672 14348 8736
rect 14412 8672 14428 8736
rect 14492 8672 14508 8736
rect 14572 8672 14580 8736
rect 14260 7648 14580 8672
rect 14260 7584 14268 7648
rect 14332 7584 14348 7648
rect 14412 7584 14428 7648
rect 14492 7584 14508 7648
rect 14572 7584 14580 7648
rect 14260 6560 14580 7584
rect 14260 6496 14268 6560
rect 14332 6496 14348 6560
rect 14412 6496 14428 6560
rect 14492 6496 14508 6560
rect 14572 6496 14580 6560
rect 14260 5472 14580 6496
rect 14260 5408 14268 5472
rect 14332 5408 14348 5472
rect 14412 5408 14428 5472
rect 14492 5408 14508 5472
rect 14572 5408 14580 5472
rect 14260 4384 14580 5408
rect 14260 4320 14268 4384
rect 14332 4320 14348 4384
rect 14412 4320 14428 4384
rect 14492 4320 14508 4384
rect 14572 4320 14580 4384
rect 14260 3296 14580 4320
rect 14260 3232 14268 3296
rect 14332 3232 14348 3296
rect 14412 3232 14428 3296
rect 14492 3232 14508 3296
rect 14572 3232 14580 3296
rect 14260 2208 14580 3232
rect 14260 2144 14268 2208
rect 14332 2144 14348 2208
rect 14412 2144 14428 2208
rect 14492 2144 14508 2208
rect 14572 2144 14580 2208
rect 14260 2128 14580 2144
rect 16480 47360 16800 47376
rect 16480 47296 16488 47360
rect 16552 47296 16568 47360
rect 16632 47296 16648 47360
rect 16712 47296 16728 47360
rect 16792 47296 16800 47360
rect 16480 46272 16800 47296
rect 16480 46208 16488 46272
rect 16552 46208 16568 46272
rect 16632 46208 16648 46272
rect 16712 46208 16728 46272
rect 16792 46208 16800 46272
rect 16480 45184 16800 46208
rect 16480 45120 16488 45184
rect 16552 45120 16568 45184
rect 16632 45120 16648 45184
rect 16712 45120 16728 45184
rect 16792 45120 16800 45184
rect 16480 44096 16800 45120
rect 16480 44032 16488 44096
rect 16552 44032 16568 44096
rect 16632 44032 16648 44096
rect 16712 44032 16728 44096
rect 16792 44032 16800 44096
rect 16480 43008 16800 44032
rect 16480 42944 16488 43008
rect 16552 42944 16568 43008
rect 16632 42944 16648 43008
rect 16712 42944 16728 43008
rect 16792 42944 16800 43008
rect 16480 41920 16800 42944
rect 16480 41856 16488 41920
rect 16552 41856 16568 41920
rect 16632 41856 16648 41920
rect 16712 41856 16728 41920
rect 16792 41856 16800 41920
rect 16480 40832 16800 41856
rect 16480 40768 16488 40832
rect 16552 40768 16568 40832
rect 16632 40768 16648 40832
rect 16712 40768 16728 40832
rect 16792 40768 16800 40832
rect 16480 39744 16800 40768
rect 16480 39680 16488 39744
rect 16552 39680 16568 39744
rect 16632 39680 16648 39744
rect 16712 39680 16728 39744
rect 16792 39680 16800 39744
rect 16480 38656 16800 39680
rect 16480 38592 16488 38656
rect 16552 38592 16568 38656
rect 16632 38592 16648 38656
rect 16712 38592 16728 38656
rect 16792 38592 16800 38656
rect 16480 37568 16800 38592
rect 16480 37504 16488 37568
rect 16552 37504 16568 37568
rect 16632 37504 16648 37568
rect 16712 37504 16728 37568
rect 16792 37504 16800 37568
rect 16480 36480 16800 37504
rect 16480 36416 16488 36480
rect 16552 36416 16568 36480
rect 16632 36416 16648 36480
rect 16712 36416 16728 36480
rect 16792 36416 16800 36480
rect 16480 35392 16800 36416
rect 16480 35328 16488 35392
rect 16552 35328 16568 35392
rect 16632 35328 16648 35392
rect 16712 35328 16728 35392
rect 16792 35328 16800 35392
rect 16480 34304 16800 35328
rect 16480 34240 16488 34304
rect 16552 34240 16568 34304
rect 16632 34240 16648 34304
rect 16712 34240 16728 34304
rect 16792 34240 16800 34304
rect 16480 33216 16800 34240
rect 16480 33152 16488 33216
rect 16552 33152 16568 33216
rect 16632 33152 16648 33216
rect 16712 33152 16728 33216
rect 16792 33152 16800 33216
rect 16480 32128 16800 33152
rect 16480 32064 16488 32128
rect 16552 32064 16568 32128
rect 16632 32064 16648 32128
rect 16712 32064 16728 32128
rect 16792 32064 16800 32128
rect 16480 31040 16800 32064
rect 16480 30976 16488 31040
rect 16552 30976 16568 31040
rect 16632 30976 16648 31040
rect 16712 30976 16728 31040
rect 16792 30976 16800 31040
rect 16480 29952 16800 30976
rect 16480 29888 16488 29952
rect 16552 29888 16568 29952
rect 16632 29888 16648 29952
rect 16712 29888 16728 29952
rect 16792 29888 16800 29952
rect 16480 28864 16800 29888
rect 16480 28800 16488 28864
rect 16552 28800 16568 28864
rect 16632 28800 16648 28864
rect 16712 28800 16728 28864
rect 16792 28800 16800 28864
rect 16480 27776 16800 28800
rect 16480 27712 16488 27776
rect 16552 27712 16568 27776
rect 16632 27712 16648 27776
rect 16712 27712 16728 27776
rect 16792 27712 16800 27776
rect 16480 26688 16800 27712
rect 16480 26624 16488 26688
rect 16552 26624 16568 26688
rect 16632 26624 16648 26688
rect 16712 26624 16728 26688
rect 16792 26624 16800 26688
rect 16480 25600 16800 26624
rect 16480 25536 16488 25600
rect 16552 25536 16568 25600
rect 16632 25536 16648 25600
rect 16712 25536 16728 25600
rect 16792 25536 16800 25600
rect 16480 24512 16800 25536
rect 16480 24448 16488 24512
rect 16552 24448 16568 24512
rect 16632 24448 16648 24512
rect 16712 24448 16728 24512
rect 16792 24448 16800 24512
rect 16480 23424 16800 24448
rect 16480 23360 16488 23424
rect 16552 23360 16568 23424
rect 16632 23360 16648 23424
rect 16712 23360 16728 23424
rect 16792 23360 16800 23424
rect 16480 22336 16800 23360
rect 16480 22272 16488 22336
rect 16552 22272 16568 22336
rect 16632 22272 16648 22336
rect 16712 22272 16728 22336
rect 16792 22272 16800 22336
rect 16480 21248 16800 22272
rect 16480 21184 16488 21248
rect 16552 21184 16568 21248
rect 16632 21184 16648 21248
rect 16712 21184 16728 21248
rect 16792 21184 16800 21248
rect 16480 20160 16800 21184
rect 16480 20096 16488 20160
rect 16552 20096 16568 20160
rect 16632 20096 16648 20160
rect 16712 20096 16728 20160
rect 16792 20096 16800 20160
rect 16480 19072 16800 20096
rect 16480 19008 16488 19072
rect 16552 19008 16568 19072
rect 16632 19008 16648 19072
rect 16712 19008 16728 19072
rect 16792 19008 16800 19072
rect 16480 17984 16800 19008
rect 16480 17920 16488 17984
rect 16552 17920 16568 17984
rect 16632 17920 16648 17984
rect 16712 17920 16728 17984
rect 16792 17920 16800 17984
rect 16480 16896 16800 17920
rect 16480 16832 16488 16896
rect 16552 16832 16568 16896
rect 16632 16832 16648 16896
rect 16712 16832 16728 16896
rect 16792 16832 16800 16896
rect 16480 15808 16800 16832
rect 16480 15744 16488 15808
rect 16552 15744 16568 15808
rect 16632 15744 16648 15808
rect 16712 15744 16728 15808
rect 16792 15744 16800 15808
rect 16480 14720 16800 15744
rect 16480 14656 16488 14720
rect 16552 14656 16568 14720
rect 16632 14656 16648 14720
rect 16712 14656 16728 14720
rect 16792 14656 16800 14720
rect 16480 13632 16800 14656
rect 16480 13568 16488 13632
rect 16552 13568 16568 13632
rect 16632 13568 16648 13632
rect 16712 13568 16728 13632
rect 16792 13568 16800 13632
rect 16480 12544 16800 13568
rect 16480 12480 16488 12544
rect 16552 12480 16568 12544
rect 16632 12480 16648 12544
rect 16712 12480 16728 12544
rect 16792 12480 16800 12544
rect 16480 11456 16800 12480
rect 16480 11392 16488 11456
rect 16552 11392 16568 11456
rect 16632 11392 16648 11456
rect 16712 11392 16728 11456
rect 16792 11392 16800 11456
rect 16480 10368 16800 11392
rect 16480 10304 16488 10368
rect 16552 10304 16568 10368
rect 16632 10304 16648 10368
rect 16712 10304 16728 10368
rect 16792 10304 16800 10368
rect 16480 9280 16800 10304
rect 16480 9216 16488 9280
rect 16552 9216 16568 9280
rect 16632 9216 16648 9280
rect 16712 9216 16728 9280
rect 16792 9216 16800 9280
rect 16480 8192 16800 9216
rect 16480 8128 16488 8192
rect 16552 8128 16568 8192
rect 16632 8128 16648 8192
rect 16712 8128 16728 8192
rect 16792 8128 16800 8192
rect 16480 7104 16800 8128
rect 16480 7040 16488 7104
rect 16552 7040 16568 7104
rect 16632 7040 16648 7104
rect 16712 7040 16728 7104
rect 16792 7040 16800 7104
rect 16480 6016 16800 7040
rect 16480 5952 16488 6016
rect 16552 5952 16568 6016
rect 16632 5952 16648 6016
rect 16712 5952 16728 6016
rect 16792 5952 16800 6016
rect 16480 4928 16800 5952
rect 16480 4864 16488 4928
rect 16552 4864 16568 4928
rect 16632 4864 16648 4928
rect 16712 4864 16728 4928
rect 16792 4864 16800 4928
rect 16480 3840 16800 4864
rect 16480 3776 16488 3840
rect 16552 3776 16568 3840
rect 16632 3776 16648 3840
rect 16712 3776 16728 3840
rect 16792 3776 16800 3840
rect 16480 2752 16800 3776
rect 16480 2688 16488 2752
rect 16552 2688 16568 2752
rect 16632 2688 16648 2752
rect 16712 2688 16728 2752
rect 16792 2688 16800 2752
rect 16480 2128 16800 2688
rect 18699 46816 19019 47376
rect 18699 46752 18707 46816
rect 18771 46752 18787 46816
rect 18851 46752 18867 46816
rect 18931 46752 18947 46816
rect 19011 46752 19019 46816
rect 18699 45728 19019 46752
rect 18699 45664 18707 45728
rect 18771 45664 18787 45728
rect 18851 45664 18867 45728
rect 18931 45664 18947 45728
rect 19011 45664 19019 45728
rect 18699 44640 19019 45664
rect 18699 44576 18707 44640
rect 18771 44576 18787 44640
rect 18851 44576 18867 44640
rect 18931 44576 18947 44640
rect 19011 44576 19019 44640
rect 18699 43552 19019 44576
rect 18699 43488 18707 43552
rect 18771 43488 18787 43552
rect 18851 43488 18867 43552
rect 18931 43488 18947 43552
rect 19011 43488 19019 43552
rect 18699 42464 19019 43488
rect 18699 42400 18707 42464
rect 18771 42400 18787 42464
rect 18851 42400 18867 42464
rect 18931 42400 18947 42464
rect 19011 42400 19019 42464
rect 18699 41376 19019 42400
rect 18699 41312 18707 41376
rect 18771 41312 18787 41376
rect 18851 41312 18867 41376
rect 18931 41312 18947 41376
rect 19011 41312 19019 41376
rect 18699 40288 19019 41312
rect 18699 40224 18707 40288
rect 18771 40224 18787 40288
rect 18851 40224 18867 40288
rect 18931 40224 18947 40288
rect 19011 40224 19019 40288
rect 18699 39200 19019 40224
rect 18699 39136 18707 39200
rect 18771 39136 18787 39200
rect 18851 39136 18867 39200
rect 18931 39136 18947 39200
rect 19011 39136 19019 39200
rect 18699 38112 19019 39136
rect 18699 38048 18707 38112
rect 18771 38048 18787 38112
rect 18851 38048 18867 38112
rect 18931 38048 18947 38112
rect 19011 38048 19019 38112
rect 18699 37024 19019 38048
rect 18699 36960 18707 37024
rect 18771 36960 18787 37024
rect 18851 36960 18867 37024
rect 18931 36960 18947 37024
rect 19011 36960 19019 37024
rect 18699 35936 19019 36960
rect 18699 35872 18707 35936
rect 18771 35872 18787 35936
rect 18851 35872 18867 35936
rect 18931 35872 18947 35936
rect 19011 35872 19019 35936
rect 18699 34848 19019 35872
rect 18699 34784 18707 34848
rect 18771 34784 18787 34848
rect 18851 34784 18867 34848
rect 18931 34784 18947 34848
rect 19011 34784 19019 34848
rect 18699 33760 19019 34784
rect 18699 33696 18707 33760
rect 18771 33696 18787 33760
rect 18851 33696 18867 33760
rect 18931 33696 18947 33760
rect 19011 33696 19019 33760
rect 18699 32672 19019 33696
rect 18699 32608 18707 32672
rect 18771 32608 18787 32672
rect 18851 32608 18867 32672
rect 18931 32608 18947 32672
rect 19011 32608 19019 32672
rect 18699 31584 19019 32608
rect 18699 31520 18707 31584
rect 18771 31520 18787 31584
rect 18851 31520 18867 31584
rect 18931 31520 18947 31584
rect 19011 31520 19019 31584
rect 18699 30496 19019 31520
rect 18699 30432 18707 30496
rect 18771 30432 18787 30496
rect 18851 30432 18867 30496
rect 18931 30432 18947 30496
rect 19011 30432 19019 30496
rect 18699 29408 19019 30432
rect 18699 29344 18707 29408
rect 18771 29344 18787 29408
rect 18851 29344 18867 29408
rect 18931 29344 18947 29408
rect 19011 29344 19019 29408
rect 18699 28320 19019 29344
rect 18699 28256 18707 28320
rect 18771 28256 18787 28320
rect 18851 28256 18867 28320
rect 18931 28256 18947 28320
rect 19011 28256 19019 28320
rect 18699 27232 19019 28256
rect 18699 27168 18707 27232
rect 18771 27168 18787 27232
rect 18851 27168 18867 27232
rect 18931 27168 18947 27232
rect 19011 27168 19019 27232
rect 18699 26144 19019 27168
rect 18699 26080 18707 26144
rect 18771 26080 18787 26144
rect 18851 26080 18867 26144
rect 18931 26080 18947 26144
rect 19011 26080 19019 26144
rect 18699 25056 19019 26080
rect 18699 24992 18707 25056
rect 18771 24992 18787 25056
rect 18851 24992 18867 25056
rect 18931 24992 18947 25056
rect 19011 24992 19019 25056
rect 18699 23968 19019 24992
rect 18699 23904 18707 23968
rect 18771 23904 18787 23968
rect 18851 23904 18867 23968
rect 18931 23904 18947 23968
rect 19011 23904 19019 23968
rect 18699 22880 19019 23904
rect 18699 22816 18707 22880
rect 18771 22816 18787 22880
rect 18851 22816 18867 22880
rect 18931 22816 18947 22880
rect 19011 22816 19019 22880
rect 18699 21792 19019 22816
rect 18699 21728 18707 21792
rect 18771 21728 18787 21792
rect 18851 21728 18867 21792
rect 18931 21728 18947 21792
rect 19011 21728 19019 21792
rect 18699 20704 19019 21728
rect 18699 20640 18707 20704
rect 18771 20640 18787 20704
rect 18851 20640 18867 20704
rect 18931 20640 18947 20704
rect 19011 20640 19019 20704
rect 18699 19616 19019 20640
rect 18699 19552 18707 19616
rect 18771 19552 18787 19616
rect 18851 19552 18867 19616
rect 18931 19552 18947 19616
rect 19011 19552 19019 19616
rect 18699 18528 19019 19552
rect 18699 18464 18707 18528
rect 18771 18464 18787 18528
rect 18851 18464 18867 18528
rect 18931 18464 18947 18528
rect 19011 18464 19019 18528
rect 18699 17440 19019 18464
rect 18699 17376 18707 17440
rect 18771 17376 18787 17440
rect 18851 17376 18867 17440
rect 18931 17376 18947 17440
rect 19011 17376 19019 17440
rect 18699 16352 19019 17376
rect 18699 16288 18707 16352
rect 18771 16288 18787 16352
rect 18851 16288 18867 16352
rect 18931 16288 18947 16352
rect 19011 16288 19019 16352
rect 18699 15264 19019 16288
rect 18699 15200 18707 15264
rect 18771 15200 18787 15264
rect 18851 15200 18867 15264
rect 18931 15200 18947 15264
rect 19011 15200 19019 15264
rect 18699 14176 19019 15200
rect 18699 14112 18707 14176
rect 18771 14112 18787 14176
rect 18851 14112 18867 14176
rect 18931 14112 18947 14176
rect 19011 14112 19019 14176
rect 18699 13088 19019 14112
rect 18699 13024 18707 13088
rect 18771 13024 18787 13088
rect 18851 13024 18867 13088
rect 18931 13024 18947 13088
rect 19011 13024 19019 13088
rect 18699 12000 19019 13024
rect 18699 11936 18707 12000
rect 18771 11936 18787 12000
rect 18851 11936 18867 12000
rect 18931 11936 18947 12000
rect 19011 11936 19019 12000
rect 18699 10912 19019 11936
rect 18699 10848 18707 10912
rect 18771 10848 18787 10912
rect 18851 10848 18867 10912
rect 18931 10848 18947 10912
rect 19011 10848 19019 10912
rect 18699 9824 19019 10848
rect 18699 9760 18707 9824
rect 18771 9760 18787 9824
rect 18851 9760 18867 9824
rect 18931 9760 18947 9824
rect 19011 9760 19019 9824
rect 18699 8736 19019 9760
rect 18699 8672 18707 8736
rect 18771 8672 18787 8736
rect 18851 8672 18867 8736
rect 18931 8672 18947 8736
rect 19011 8672 19019 8736
rect 18699 7648 19019 8672
rect 18699 7584 18707 7648
rect 18771 7584 18787 7648
rect 18851 7584 18867 7648
rect 18931 7584 18947 7648
rect 19011 7584 19019 7648
rect 18699 6560 19019 7584
rect 18699 6496 18707 6560
rect 18771 6496 18787 6560
rect 18851 6496 18867 6560
rect 18931 6496 18947 6560
rect 19011 6496 19019 6560
rect 18699 5472 19019 6496
rect 18699 5408 18707 5472
rect 18771 5408 18787 5472
rect 18851 5408 18867 5472
rect 18931 5408 18947 5472
rect 19011 5408 19019 5472
rect 18699 4384 19019 5408
rect 18699 4320 18707 4384
rect 18771 4320 18787 4384
rect 18851 4320 18867 4384
rect 18931 4320 18947 4384
rect 19011 4320 19019 4384
rect 18699 3296 19019 4320
rect 18699 3232 18707 3296
rect 18771 3232 18787 3296
rect 18851 3232 18867 3296
rect 18931 3232 18947 3296
rect 19011 3232 19019 3296
rect 18699 2208 19019 3232
rect 18699 2144 18707 2208
rect 18771 2144 18787 2208
rect 18851 2144 18867 2208
rect 18931 2144 18947 2208
rect 19011 2144 19019 2208
rect 18699 2128 19019 2144
use sky130_fd_sc_hd__nor2_1  _09_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _10_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _11_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _12_
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _13_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16376 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _14_
timestamp 1688980957
transform -1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_1  _15_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17848 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _16_
timestamp 1688980957
transform 1 0 17664 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _17_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_1  _18_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _19_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15732 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _20_
timestamp 1688980957
transform -1 0 16376 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _21_
timestamp 1688980957
transform 1 0 16928 0 -1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold2_A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold6_A
timestamp 1688980957
transform -1 0 18584 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output4_A
timestamp 1688980957
transform -1 0 17112 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_A
timestamp 1688980957
transform -1 0 18584 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1688980957
transform -1 0 17480 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1688980957
transform -1 0 17480 0 1 5440
box -38 -48 1878 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 1688980957
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_149 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_154
timestamp 1688980957
transform 1 0 15272 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1688980957
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_185
timestamp 1688980957
transform 1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_173
timestamp 1688980957
transform 1 0 17020 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_186
timestamp 1688980957
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_178
timestamp 1688980957
transform 1 0 17480 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_189
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_187
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 1688980957
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_157
timestamp 1688980957
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_163
timestamp 1688980957
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_187
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_189
timestamp 1688980957
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 1688980957
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1688980957
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_189
timestamp 1688980957
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 1688980957
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 1688980957
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 1688980957
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 1688980957
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_189
timestamp 1688980957
transform 1 0 18492 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 1688980957
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 1688980957
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_173
timestamp 1688980957
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 1688980957
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 1688980957
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1688980957
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 1688980957
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 1688980957
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 1688980957
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 1688980957
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_189
timestamp 1688980957
transform 1 0 18492 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 1688980957
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1688980957
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1688980957
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1688980957
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 1688980957
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 1688980957
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_189
timestamp 1688980957
transform 1 0 18492 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 1688980957
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 1688980957
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 1688980957
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 1688980957
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_189
timestamp 1688980957
transform 1 0 18492 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 1688980957
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 1688980957
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 1688980957
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 1688980957
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 1688980957
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 1688980957
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 1688980957
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_189
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 1688980957
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 1688980957
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 1688980957
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 1688980957
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 1688980957
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_189
timestamp 1688980957
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 1688980957
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 1688980957
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 1688980957
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_189
timestamp 1688980957
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 1688980957
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 1688980957
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 1688980957
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_185
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 1688980957
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 1688980957
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_189
timestamp 1688980957
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 1688980957
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 1688980957
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 1688980957
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 1688980957
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 1688980957
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_189
timestamp 1688980957
transform 1 0 18492 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 1688980957
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_189
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 1688980957
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 1688980957
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 1688980957
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_189
timestamp 1688980957
transform 1 0 18492 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 1688980957
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 1688980957
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_189
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 1688980957
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 1688980957
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 1688980957
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 1688980957
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 1688980957
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 1688980957
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_189
timestamp 1688980957
transform 1 0 18492 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 1688980957
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 1688980957
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 1688980957
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 1688980957
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 1688980957
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_189
timestamp 1688980957
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 1688980957
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 1688980957
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 1688980957
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_189
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 1688980957
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 1688980957
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 1688980957
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_171
timestamp 1688980957
transform 1 0 16836 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 1688980957
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_189
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 1688980957
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 1688980957
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 1688980957
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 1688980957
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 1688980957
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 1688980957
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 1688980957
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 1688980957
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_189
timestamp 1688980957
transform 1 0 18492 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 1688980957
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 1688980957
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 1688980957
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_189
timestamp 1688980957
transform 1 0 18492 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_189
timestamp 1688980957
transform 1 0 18492 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_189
timestamp 1688980957
transform 1 0 18492 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 1688980957
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 1688980957
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 1688980957
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 1688980957
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_189
timestamp 1688980957
transform 1 0 18492 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_189
timestamp 1688980957
transform 1 0 18492 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_121
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_133
timestamp 1688980957
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_189
timestamp 1688980957
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_189
timestamp 1688980957
transform 1 0 18492 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_15
timestamp 1688980957
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_189
timestamp 1688980957
transform 1 0 18492 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_185
timestamp 1688980957
transform 1 0 18124 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_15
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_173
timestamp 1688980957
transform 1 0 17020 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_189
timestamp 1688980957
transform 1 0 18492 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_189
timestamp 1688980957
transform 1 0 18492 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_181
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_189
timestamp 1688980957
transform 1 0 18492 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1688980957
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1688980957
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1688980957
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1688980957
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1688980957
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1688980957
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1688980957
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_189
timestamp 1688980957
transform 1 0 18492 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_27
timestamp 1688980957
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_39
timestamp 1688980957
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_51
timestamp 1688980957
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1688980957
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1688980957
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1688980957
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1688980957
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_77_181
timestamp 1688980957
transform 1 0 17756 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_189
timestamp 1688980957
transform 1 0 18492 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1688980957
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1688980957
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1688980957
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1688980957
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1688980957
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1688980957
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_189
timestamp 1688980957
transform 1 0 18492 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1688980957
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1688980957
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1688980957
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 1688980957
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 1688980957
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1688980957
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1688980957
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1688980957
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_181
timestamp 1688980957
transform 1 0 17756 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_189
timestamp 1688980957
transform 1 0 18492 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_3
timestamp 1688980957
transform 1 0 1380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_15
timestamp 1688980957
transform 1 0 2484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1688980957
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1688980957
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1688980957
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1688980957
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1688980957
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1688980957
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1688980957
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1688980957
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1688980957
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1688980957
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1688980957
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1688980957
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_189
timestamp 1688980957
transform 1 0 18492 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1688980957
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1688980957
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1688980957
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1688980957
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 1688980957
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1688980957
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1688980957
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1688980957
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1688980957
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1688980957
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1688980957
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1688980957
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1688980957
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1688980957
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1688980957
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1688980957
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1688980957
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1688980957
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1688980957
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_81_181
timestamp 1688980957
transform 1 0 17756 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_189
timestamp 1688980957
transform 1 0 18492 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1688980957
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1688980957
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1688980957
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1688980957
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1688980957
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_53
timestamp 1688980957
transform 1 0 5980 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_57
timestamp 1688980957
transform 1 0 6348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_69
timestamp 1688980957
transform 1 0 7452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_81
timestamp 1688980957
transform 1 0 8556 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1688980957
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1688980957
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_109
timestamp 1688980957
transform 1 0 11132 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_113
timestamp 1688980957
transform 1 0 11500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_125
timestamp 1688980957
transform 1 0 12604 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_137
timestamp 1688980957
transform 1 0 13708 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1688980957
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1688980957
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_82_165
timestamp 1688980957
transform 1 0 16284 0 1 46784
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_169
timestamp 1688980957
transform 1 0 16652 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_181
timestamp 1688980957
transform 1 0 17756 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  hold2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16376 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 16836 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 18584 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 17848 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform -1 0 18216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1688980957
transform 1 0 14996 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17112 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output3
timestamp 1688980957
transform 1 0 17112 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output4
timestamp 1688980957
transform 1 0 17112 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output5
timestamp 1688980957
transform -1 0 18584 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 18860 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 18860 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 18860 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 18860 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 18860 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 18860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 18860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 18860 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 18860 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 18860 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 18860 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 18860 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 18860 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 18860 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 18860 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 18860 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 18860 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 18860 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 18860 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 18860 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 18860 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 18860 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 18860 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 18860 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 18860 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1688980957
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1688980957
transform -1 0 18860 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1688980957
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1688980957
transform -1 0 18860 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  user_proj_example_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  user_proj_example_7
timestamp 1688980957
transform 1 0 18308 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  user_proj_example_8
timestamp 1688980957
transform 1 0 18308 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  user_proj_example_9
timestamp 1688980957
transform 1 0 18308 0 1 46784
box -38 -48 314 592
<< labels >>
flabel metal3 s 19200 9256 20000 9376 0 FreeSans 480 0 0 0 io_oeb[0]
port 0 nsew signal tristate
flabel metal3 s 19200 21768 20000 21888 0 FreeSans 480 0 0 0 io_oeb[1]
port 1 nsew signal tristate
flabel metal3 s 19200 34280 20000 34400 0 FreeSans 480 0 0 0 io_oeb[2]
port 2 nsew signal tristate
flabel metal3 s 19200 46792 20000 46912 0 FreeSans 480 0 0 0 io_oeb[3]
port 3 nsew signal tristate
flabel metal3 s 19200 3000 20000 3120 0 FreeSans 480 0 0 0 io_out[0]
port 4 nsew signal tristate
flabel metal3 s 19200 15512 20000 15632 0 FreeSans 480 0 0 0 io_out[1]
port 5 nsew signal tristate
flabel metal3 s 19200 28024 20000 28144 0 FreeSans 480 0 0 0 io_out[2]
port 6 nsew signal tristate
flabel metal3 s 19200 40536 20000 40656 0 FreeSans 480 0 0 0 io_out[3]
port 7 nsew signal tristate
flabel metal4 s 3163 2128 3483 47376 0 FreeSans 1920 90 0 0 vccd1
port 8 nsew power bidirectional
flabel metal4 s 7602 2128 7922 47376 0 FreeSans 1920 90 0 0 vccd1
port 8 nsew power bidirectional
flabel metal4 s 12041 2128 12361 47376 0 FreeSans 1920 90 0 0 vccd1
port 8 nsew power bidirectional
flabel metal4 s 16480 2128 16800 47376 0 FreeSans 1920 90 0 0 vccd1
port 8 nsew power bidirectional
flabel metal4 s 5382 2128 5702 47376 0 FreeSans 1920 90 0 0 vssd1
port 9 nsew ground bidirectional
flabel metal4 s 9821 2128 10141 47376 0 FreeSans 1920 90 0 0 vssd1
port 9 nsew ground bidirectional
flabel metal4 s 14260 2128 14580 47376 0 FreeSans 1920 90 0 0 vssd1
port 9 nsew ground bidirectional
flabel metal4 s 18699 2128 19019 47376 0 FreeSans 1920 90 0 0 vssd1
port 9 nsew ground bidirectional
flabel metal2 s 4986 0 5042 800 0 FreeSans 224 90 0 0 wb_clk_i
port 10 nsew signal input
flabel metal2 s 14922 0 14978 800 0 FreeSans 224 90 0 0 wb_rst_i
port 11 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 50000
<< end >>
